`timescale 1ns / 1ps

module fi_address(
    input [15:0] angle,
    input valid_point,
    
    output [11:0] address
);
    
wire [2081:0] fi_addres;    

encoder #(
    .LEN_IN(2082)) encoder_fi_address (
    .in(fi_addres),
    .out(address)
);
    
assign fi_addres[0] = valid_point & (angle >= 16'd0 & angle <= 16'd1);
assign fi_addres[1] = valid_point & (angle > 16'd1 & angle <= 16'd23);
assign fi_addres[2] = valid_point & (angle > 16'd23 & angle <= 16'd40);
assign fi_addres[3] = valid_point & (angle > 16'd40 & angle <= 16'd56);
assign fi_addres[4] = valid_point & (angle > 16'd56 & angle <= 16'd77);
assign fi_addres[5] = valid_point & (angle > 16'd77 & angle <= 16'd95);
assign fi_addres[6] = valid_point & (angle > 16'd95 & angle <= 16'd113);
assign fi_addres[7] = valid_point & (angle > 16'd113 & angle <= 16'd137);
assign fi_addres[8] = valid_point & (angle > 16'd137 & angle <= 16'd155);
assign fi_addres[9] = valid_point & (angle > 16'd155 & angle <= 16'd173);
assign fi_addres[10] = valid_point & (angle > 16'd173 & angle <= 16'd191);
assign fi_addres[11] = valid_point & (angle > 16'd191 & angle <= 16'd208);
assign fi_addres[12] = valid_point & (angle > 16'd208 & angle <= 16'd226);
assign fi_addres[13] = valid_point & (angle > 16'd226 & angle <= 16'd258);
assign fi_addres[14] = valid_point & (angle > 16'd258 & angle <= 16'd276);
assign fi_addres[15] = valid_point & (angle > 16'd276 & angle <= 16'd307);
assign fi_addres[16] = valid_point & (angle > 16'd307 & angle <= 16'd326);
assign fi_addres[17] = valid_point & (angle > 16'd326 & angle <= 16'd344);
assign fi_addres[18] = valid_point & (angle > 16'd344 & angle <= 16'd362);
assign fi_addres[19] = valid_point & (angle > 16'd362 & angle <= 16'd389);
assign fi_addres[20] = valid_point & (angle > 16'd389 & angle <= 16'd407);
assign fi_addres[21] = valid_point & (angle > 16'd407 & angle <= 16'd424);
assign fi_addres[22] = valid_point & (angle > 16'd424 & angle <= 16'd456);
assign fi_addres[23] = valid_point & (angle > 16'd456 & angle <= 16'd474);
assign fi_addres[24] = valid_point & (angle > 16'd474 & angle <= 16'd492);
assign fi_addres[25] = valid_point & (angle > 16'd492 & angle <= 16'd524);
assign fi_addres[26] = valid_point & (angle > 16'd524 & angle <= 16'd542);
assign fi_addres[27] = valid_point & (angle > 16'd542 & angle <= 16'd560);
assign fi_addres[28] = valid_point & (angle > 16'd560 & angle <= 16'd578);
assign fi_addres[29] = valid_point & (angle > 16'd578 & angle <= 16'd596);
assign fi_addres[30] = valid_point & (angle > 16'd596 & angle <= 16'd623);
assign fi_addres[31] = valid_point & (angle > 16'd623 & angle <= 16'd640);
assign fi_addres[32] = valid_point & (angle > 16'd640 & angle <= 16'd659);
assign fi_addres[33] = valid_point & (angle > 16'd659 & angle <= 16'd677);
assign fi_addres[34] = valid_point & (angle > 16'd677 & angle <= 16'd695);
assign fi_addres[35] = valid_point & (angle > 16'd695 & angle <= 16'd716);
assign fi_addres[36] = valid_point & (angle > 16'd716 & angle <= 16'd745);
assign fi_addres[37] = valid_point & (angle > 16'd745 & angle <= 16'd762);
assign fi_addres[38] = valid_point & (angle > 16'd762 & angle <= 16'd788);
assign fi_addres[39] = valid_point & (angle > 16'd788 & angle <= 16'd804);
assign fi_addres[40] = valid_point & (angle > 16'd804 & angle <= 16'd822);
assign fi_addres[41] = valid_point & (angle > 16'd822 & angle <= 16'd840);
assign fi_addres[42] = valid_point & (angle > 16'd840 & angle <= 16'd858);
assign fi_addres[43] = valid_point & (angle > 16'd858 & angle <= 16'd876);
assign fi_addres[44] = valid_point & (angle > 16'd876 & angle <= 16'd894);
assign fi_addres[45] = valid_point & (angle > 16'd894 & angle <= 16'd903);
assign fi_addres[46] = valid_point & (angle > 16'd903 & angle <= 16'd921);
assign fi_addres[47] = valid_point & (angle > 16'd921 & angle <= 16'd939);
assign fi_addres[48] = valid_point & (angle > 16'd939 & angle <= 16'd957);
assign fi_addres[49] = valid_point & (angle > 16'd957 & angle <= 16'd975);
assign fi_addres[50] = valid_point & (angle > 16'd975 & angle <= 16'd993);
assign fi_addres[51] = valid_point & (angle > 16'd993 & angle <= 16'd1011);
assign fi_addres[52] = valid_point & (angle > 16'd1011 & angle <= 16'd1020);
assign fi_addres[53] = valid_point & (angle > 16'd1020 & angle <= 16'd1038);
assign fi_addres[54] = valid_point & (angle > 16'd1038 & angle <= 16'd1068);
assign fi_addres[55] = valid_point & (angle > 16'd1068 & angle <= 16'd1092);
assign fi_addres[56] = valid_point & (angle > 16'd1092 & angle <= 16'd1110);
assign fi_addres[57] = valid_point & (angle > 16'd1110 & angle <= 16'd1128);
assign fi_addres[58] = valid_point & (angle > 16'd1128 & angle <= 16'd1137);
assign fi_addres[59] = valid_point & (angle > 16'd1137 & angle <= 16'd1155);
assign fi_addres[60] = valid_point & (angle > 16'd1155 & angle <= 16'd1173);
assign fi_addres[61] = valid_point & (angle > 16'd1173 & angle <= 16'd1191);
assign fi_addres[62] = valid_point & (angle > 16'd1191 & angle <= 16'd1209);
assign fi_addres[63] = valid_point & (angle > 16'd1209 & angle <= 16'd1227);
assign fi_addres[64] = valid_point & (angle > 16'd1227 & angle <= 16'd1245);
assign fi_addres[65] = valid_point & (angle > 16'd1245 & angle <= 16'd1254);
assign fi_addres[66] = valid_point & (angle > 16'd1254 & angle <= 16'd1272);
assign fi_addres[67] = valid_point & (angle > 16'd1272 & angle <= 16'd1290);
assign fi_addres[68] = valid_point & (angle > 16'd1290 & angle <= 16'd1308);
assign fi_addres[69] = valid_point & (angle > 16'd1308 & angle <= 16'd1326);
assign fi_addres[70] = valid_point & (angle > 16'd1326 & angle <= 16'd1344);
assign fi_addres[71] = valid_point & (angle > 16'd1344 & angle <= 16'd1362);
assign fi_addres[72] = valid_point & (angle > 16'd1362 & angle <= 16'd1380);
assign fi_addres[73] = valid_point & (angle > 16'd1380 & angle <= 16'd1389);
assign fi_addres[74] = valid_point & (angle > 16'd1389 & angle <= 16'd1407);
assign fi_addres[75] = valid_point & (angle > 16'd1407 & angle <= 16'd1425);
assign fi_addres[76] = valid_point & (angle > 16'd1425 & angle <= 16'd1443);
assign fi_addres[77] = valid_point & (angle > 16'd1443 & angle <= 16'd1460);
assign fi_addres[78] = valid_point & (angle > 16'd1460 & angle <= 16'd1478);
assign fi_addres[79] = valid_point & (angle > 16'd1478 & angle <= 16'd1496);
assign fi_addres[80] = valid_point & (angle > 16'd1496 & angle <= 16'd1505);
assign fi_addres[81] = valid_point & (angle > 16'd1505 & angle <= 16'd1523);
assign fi_addres[82] = valid_point & (angle > 16'd1523 & angle <= 16'd1541);
assign fi_addres[83] = valid_point & (angle > 16'd1541 & angle <= 16'd1559);
assign fi_addres[84] = valid_point & (angle > 16'd1559 & angle <= 16'd1577);
assign fi_addres[85] = valid_point & (angle > 16'd1577 & angle <= 16'd1595);
assign fi_addres[86] = valid_point & (angle > 16'd1595 & angle <= 16'd1613);
assign fi_addres[87] = valid_point & (angle > 16'd1613 & angle <= 16'd1622);
assign fi_addres[88] = valid_point & (angle > 16'd1622 & angle <= 16'd1640);
assign fi_addres[89] = valid_point & (angle > 16'd1640 & angle <= 16'd1658);
assign fi_addres[90] = valid_point & (angle > 16'd1658 & angle <= 16'd1676);
assign fi_addres[91] = valid_point & (angle > 16'd1676 & angle <= 16'd1694);
assign fi_addres[92] = valid_point & (angle > 16'd1694 & angle <= 16'd1712);
assign fi_addres[93] = valid_point & (angle > 16'd1712 & angle <= 16'd1730);
assign fi_addres[94] = valid_point & (angle > 16'd1730 & angle <= 16'd1739);
assign fi_addres[95] = valid_point & (angle > 16'd1739 & angle <= 16'd1757);
assign fi_addres[96] = valid_point & (angle > 16'd1757 & angle <= 16'd1775);
assign fi_addres[97] = valid_point & (angle > 16'd1775 & angle <= 16'd1793);
assign fi_addres[98] = valid_point & (angle > 16'd1793 & angle <= 16'd1811);
assign fi_addres[99] = valid_point & (angle > 16'd1811 & angle <= 16'd1829);
assign fi_addres[100] = valid_point & (angle > 16'd1829 & angle <= 16'd1847);
assign fi_addres[101] = valid_point & (angle > 16'd1847 & angle <= 16'd1856);
assign fi_addres[102] = valid_point & (angle > 16'd1856 & angle <= 16'd1874);
assign fi_addres[103] = valid_point & (angle > 16'd1874 & angle <= 16'd1892);
assign fi_addres[104] = valid_point & (angle > 16'd1892 & angle <= 16'd1910);
assign fi_addres[105] = valid_point & (angle > 16'd1910 & angle <= 16'd1928);
assign fi_addres[106] = valid_point & (angle > 16'd1928 & angle <= 16'd1946);
assign fi_addres[107] = valid_point & (angle > 16'd1946 & angle <= 16'd1964);
assign fi_addres[108] = valid_point & (angle > 16'd1964 & angle <= 16'd1982);
assign fi_addres[109] = valid_point & (angle > 16'd1982 & angle <= 16'd1991);
assign fi_addres[110] = valid_point & (angle > 16'd1991 & angle <= 16'd2009);
assign fi_addres[111] = valid_point & (angle > 16'd2009 & angle <= 16'd2027);
assign fi_addres[112] = valid_point & (angle > 16'd2027 & angle <= 16'd2045);
assign fi_addres[113] = valid_point & (angle > 16'd2045 & angle <= 16'd2063);
assign fi_addres[114] = valid_point & (angle > 16'd2063 & angle <= 16'd2081);
assign fi_addres[115] = valid_point & (angle > 16'd2081 & angle <= 16'd2099);
assign fi_addres[116] = valid_point & (angle > 16'd2099 & angle <= 16'd2108);
assign fi_addres[117] = valid_point & (angle > 16'd2108 & angle <= 16'd2126);
assign fi_addres[118] = valid_point & (angle > 16'd2126 & angle <= 16'd2144);
assign fi_addres[119] = valid_point & (angle > 16'd2144 & angle <= 16'd2162);
assign fi_addres[120] = valid_point & (angle > 16'd2162 & angle <= 16'd2179);
assign fi_addres[121] = valid_point & (angle > 16'd2179 & angle <= 16'd2198);
assign fi_addres[122] = valid_point & (angle > 16'd2198 & angle <= 16'd2216);
assign fi_addres[123] = valid_point & (angle > 16'd2216 & angle <= 16'd2225);
assign fi_addres[124] = valid_point & (angle > 16'd2225 & angle <= 16'd2243);
assign fi_addres[125] = valid_point & (angle > 16'd2243 & angle <= 16'd2260);
assign fi_addres[126] = valid_point & (angle > 16'd2260 & angle <= 16'd2279);
assign fi_addres[127] = valid_point & (angle > 16'd2279 & angle <= 16'd2297);
assign fi_addres[128] = valid_point & (angle > 16'd2297 & angle <= 16'd2315);
assign fi_addres[129] = valid_point & (angle > 16'd2315 & angle <= 16'd2332);
assign fi_addres[130] = valid_point & (angle > 16'd2332 & angle <= 16'd2342);
assign fi_addres[131] = valid_point & (angle > 16'd2342 & angle <= 16'd2360);
assign fi_addres[132] = valid_point & (angle > 16'd2360 & angle <= 16'd2377);
assign fi_addres[133] = valid_point & (angle > 16'd2377 & angle <= 16'd2395);
assign fi_addres[134] = valid_point & (angle > 16'd2395 & angle <= 16'd2414);
assign fi_addres[135] = valid_point & (angle > 16'd2414 & angle <= 16'd2432);
assign fi_addres[136] = valid_point & (angle > 16'd2432 & angle <= 16'd2450);
assign fi_addres[137] = valid_point & (angle > 16'd2450 & angle <= 16'd2459);
assign fi_addres[138] = valid_point & (angle > 16'd2459 & angle <= 16'd2477);
assign fi_addres[139] = valid_point & (angle > 16'd2477 & angle <= 16'd2495);
assign fi_addres[140] = valid_point & (angle > 16'd2495 & angle <= 16'd2513);
assign fi_addres[141] = valid_point & (angle > 16'd2513 & angle <= 16'd2531);
assign fi_addres[142] = valid_point & (angle > 16'd2531 & angle <= 16'd2549);
assign fi_addres[143] = valid_point & (angle > 16'd2549 & angle <= 16'd2567);
assign fi_addres[144] = valid_point & (angle > 16'd2567 & angle <= 16'd2585);
assign fi_addres[145] = valid_point & (angle > 16'd2585 & angle <= 16'd2594);
assign fi_addres[146] = valid_point & (angle > 16'd2594 & angle <= 16'd2612);
assign fi_addres[147] = valid_point & (angle > 16'd2612 & angle <= 16'd2630);
assign fi_addres[148] = valid_point & (angle > 16'd2630 & angle <= 16'd2647);
assign fi_addres[149] = valid_point & (angle > 16'd2647 & angle <= 16'd2666);
assign fi_addres[150] = valid_point & (angle > 16'd2666 & angle <= 16'd2683);
assign fi_addres[151] = valid_point & (angle > 16'd2683 & angle <= 16'd2702);
assign fi_addres[152] = valid_point & (angle > 16'd2702 & angle <= 16'd2710);
assign fi_addres[153] = valid_point & (angle > 16'd2710 & angle <= 16'd2728);
assign fi_addres[154] = valid_point & (angle > 16'd2728 & angle <= 16'd2746);
assign fi_addres[155] = valid_point & (angle > 16'd2746 & angle <= 16'd2764);
assign fi_addres[156] = valid_point & (angle > 16'd2764 & angle <= 16'd2782);
assign fi_addres[157] = valid_point & (angle > 16'd2782 & angle <= 16'd2800);
assign fi_addres[158] = valid_point & (angle > 16'd2800 & angle <= 16'd2818);
assign fi_addres[159] = valid_point & (angle > 16'd2818 & angle <= 16'd2827);
assign fi_addres[160] = valid_point & (angle > 16'd2827 & angle <= 16'd2845);
assign fi_addres[161] = valid_point & (angle > 16'd2845 & angle <= 16'd2863);
assign fi_addres[162] = valid_point & (angle > 16'd2863 & angle <= 16'd2881);
assign fi_addres[163] = valid_point & (angle > 16'd2881 & angle <= 16'd2899);
assign fi_addres[164] = valid_point & (angle > 16'd2899 & angle <= 16'd2917);
assign fi_addres[165] = valid_point & (angle > 16'd2917 & angle <= 16'd2935);
assign fi_addres[166] = valid_point & (angle > 16'd2935 & angle <= 16'd2944);
assign fi_addres[167] = valid_point & (angle > 16'd2944 & angle <= 16'd2962);
assign fi_addres[168] = valid_point & (angle > 16'd2962 & angle <= 16'd2980);
assign fi_addres[169] = valid_point & (angle > 16'd2980 & angle <= 16'd2997);
assign fi_addres[170] = valid_point & (angle > 16'd2997 & angle <= 16'd3016);
assign fi_addres[171] = valid_point & (angle > 16'd3016 & angle <= 16'd3033);
assign fi_addres[172] = valid_point & (angle > 16'd3033 & angle <= 16'd3052);
assign fi_addres[173] = valid_point & (angle > 16'd3052 & angle <= 16'd3061);
assign fi_addres[174] = valid_point & (angle > 16'd3061 & angle <= 16'd3079);
assign fi_addres[175] = valid_point & (angle > 16'd3079 & angle <= 16'd3097);
assign fi_addres[176] = valid_point & (angle > 16'd3097 & angle <= 16'd3115);
assign fi_addres[177] = valid_point & (angle > 16'd3115 & angle <= 16'd3133);
assign fi_addres[178] = valid_point & (angle > 16'd3133 & angle <= 16'd3151);
assign fi_addres[179] = valid_point & (angle > 16'd3151 & angle <= 16'd3169);
assign fi_addres[180] = valid_point & (angle > 16'd3169 & angle <= 16'd3178);
assign fi_addres[181] = valid_point & (angle > 16'd3178 & angle <= 16'd3196);
assign fi_addres[182] = valid_point & (angle > 16'd3196 & angle <= 16'd3214);
assign fi_addres[183] = valid_point & (angle > 16'd3214 & angle <= 16'd3232);
assign fi_addres[184] = valid_point & (angle > 16'd3232 & angle <= 16'd3250);
assign fi_addres[185] = valid_point & (angle > 16'd3250 & angle <= 16'd3268);
assign fi_addres[186] = valid_point & (angle > 16'd3268 & angle <= 16'd3286);
assign fi_addres[187] = valid_point & (angle > 16'd3286 & angle <= 16'd3304);
assign fi_addres[188] = valid_point & (angle > 16'd3304 & angle <= 16'd3313);
assign fi_addres[189] = valid_point & (angle > 16'd3313 & angle <= 16'd3331);
assign fi_addres[190] = valid_point & (angle > 16'd3331 & angle <= 16'd3349);
assign fi_addres[191] = valid_point & (angle > 16'd3349 & angle <= 16'd3367);
assign fi_addres[192] = valid_point & (angle > 16'd3367 & angle <= 16'd3385);
assign fi_addres[193] = valid_point & (angle > 16'd3385 & angle <= 16'd3403);
assign fi_addres[194] = valid_point & (angle > 16'd3403 & angle <= 16'd3421);
assign fi_addres[195] = valid_point & (angle > 16'd3421 & angle <= 16'd3429);
assign fi_addres[196] = valid_point & (angle > 16'd3429 & angle <= 16'd3447);
assign fi_addres[197] = valid_point & (angle > 16'd3447 & angle <= 16'd3465);
assign fi_addres[198] = valid_point & (angle > 16'd3465 & angle <= 16'd3483);
assign fi_addres[199] = valid_point & (angle > 16'd3483 & angle <= 16'd3501);
assign fi_addres[200] = valid_point & (angle > 16'd3501 & angle <= 16'd3519);
assign fi_addres[201] = valid_point & (angle > 16'd3519 & angle <= 16'd3537);
assign fi_addres[202] = valid_point & (angle > 16'd3537 & angle <= 16'd3545);
assign fi_addres[203] = valid_point & (angle > 16'd3545 & angle <= 16'd3564);
assign fi_addres[204] = valid_point & (angle > 16'd3564 & angle <= 16'd3582);
assign fi_addres[205] = valid_point & (angle > 16'd3582 & angle <= 16'd3599);
assign fi_addres[206] = valid_point & (angle > 16'd3599 & angle <= 16'd3617);
assign fi_addres[207] = valid_point & (angle > 16'd3617 & angle <= 16'd3635);
assign fi_addres[208] = valid_point & (angle > 16'd3635 & angle <= 16'd3654);
assign fi_addres[209] = valid_point & (angle > 16'd3654 & angle <= 16'd3663);
assign fi_addres[210] = valid_point & (angle > 16'd3663 & angle <= 16'd3680);
assign fi_addres[211] = valid_point & (angle > 16'd3680 & angle <= 16'd3698);
assign fi_addres[212] = valid_point & (angle > 16'd3698 & angle <= 16'd3716);
assign fi_addres[213] = valid_point & (angle > 16'd3716 & angle <= 16'd3734);
assign fi_addres[214] = valid_point & (angle > 16'd3734 & angle <= 16'd3752);
assign fi_addres[215] = valid_point & (angle > 16'd3752 & angle <= 16'd3770);
assign fi_addres[216] = valid_point & (angle > 16'd3770 & angle <= 16'd3779);
assign fi_addres[217] = valid_point & (angle > 16'd3779 & angle <= 16'd3797);
assign fi_addres[218] = valid_point & (angle > 16'd3797 & angle <= 16'd3815);
assign fi_addres[219] = valid_point & (angle > 16'd3815 & angle <= 16'd3833);
assign fi_addres[220] = valid_point & (angle > 16'd3833 & angle <= 16'd3851);
assign fi_addres[221] = valid_point & (angle > 16'd3851 & angle <= 16'd3869);
assign fi_addres[222] = valid_point & (angle > 16'd3869 & angle <= 16'd3887);
assign fi_addres[223] = valid_point & (angle > 16'd3887 & angle <= 16'd3896);
assign fi_addres[224] = valid_point & (angle > 16'd3896 & angle <= 16'd3914);
assign fi_addres[225] = valid_point & (angle > 16'd3914 & angle <= 16'd3932);
assign fi_addres[226] = valid_point & (angle > 16'd3932 & angle <= 16'd3951);
assign fi_addres[227] = valid_point & (angle > 16'd3951 & angle <= 16'd3968);
assign fi_addres[228] = valid_point & (angle > 16'd3968 & angle <= 16'd3986);
assign fi_addres[229] = valid_point & (angle > 16'd3986 & angle <= 16'd4004);
assign fi_addres[230] = valid_point & (angle > 16'd4004 & angle <= 16'd4022);
assign fi_addres[231] = valid_point & (angle > 16'd4022 & angle <= 16'd4031);
assign fi_addres[232] = valid_point & (angle > 16'd4031 & angle <= 16'd4049);
assign fi_addres[233] = valid_point & (angle > 16'd4049 & angle <= 16'd4067);
assign fi_addres[234] = valid_point & (angle > 16'd4067 & angle <= 16'd4085);
assign fi_addres[235] = valid_point & (angle > 16'd4085 & angle <= 16'd4103);
assign fi_addres[236] = valid_point & (angle > 16'd4103 & angle <= 16'd4121);
assign fi_addres[237] = valid_point & (angle > 16'd4121 & angle <= 16'd4139);
assign fi_addres[238] = valid_point & (angle > 16'd4139 & angle <= 16'd4149);
assign fi_addres[239] = valid_point & (angle > 16'd4149 & angle <= 16'd4167);
assign fi_addres[240] = valid_point & (angle > 16'd4167 & angle <= 16'd4185);
assign fi_addres[241] = valid_point & (angle > 16'd4185 & angle <= 16'd4203);
assign fi_addres[242] = valid_point & (angle > 16'd4203 & angle <= 16'd4221);
assign fi_addres[243] = valid_point & (angle > 16'd4221 & angle <= 16'd4239);
assign fi_addres[244] = valid_point & (angle > 16'd4239 & angle <= 16'd4257);
assign fi_addres[245] = valid_point & (angle > 16'd4257 & angle <= 16'd4266);
assign fi_addres[246] = valid_point & (angle > 16'd4266 & angle <= 16'd4284);
assign fi_addres[247] = valid_point & (angle > 16'd4284 & angle <= 16'd4302);
assign fi_addres[248] = valid_point & (angle > 16'd4302 & angle <= 16'd4320);
assign fi_addres[249] = valid_point & (angle > 16'd4320 & angle <= 16'd4338);
assign fi_addres[250] = valid_point & (angle > 16'd4338 & angle <= 16'd4356);
assign fi_addres[251] = valid_point & (angle > 16'd4356 & angle <= 16'd4374);
assign fi_addres[252] = valid_point & (angle > 16'd4374 & angle <= 16'd4392);
assign fi_addres[253] = valid_point & (angle > 16'd4392 & angle <= 16'd4401);
assign fi_addres[254] = valid_point & (angle > 16'd4401 & angle <= 16'd4419);
assign fi_addres[255] = valid_point & (angle > 16'd4419 & angle <= 16'd4437);
assign fi_addres[256] = valid_point & (angle > 16'd4437 & angle <= 16'd4455);
assign fi_addres[257] = valid_point & (angle > 16'd4455 & angle <= 16'd4473);
assign fi_addres[258] = valid_point & (angle > 16'd4473 & angle <= 16'd4491);
assign fi_addres[259] = valid_point & (angle > 16'd4491 & angle <= 16'd4508);
assign fi_addres[260] = valid_point & (angle > 16'd4508 & angle <= 16'd4518);
assign fi_addres[261] = valid_point & (angle > 16'd4518 & angle <= 16'd4536);
assign fi_addres[262] = valid_point & (angle > 16'd4536 & angle <= 16'd4553);
assign fi_addres[263] = valid_point & (angle > 16'd4553 & angle <= 16'd4571);
assign fi_addres[264] = valid_point & (angle > 16'd4571 & angle <= 16'd4589);
assign fi_addres[265] = valid_point & (angle > 16'd4589 & angle <= 16'd4607);
assign fi_addres[266] = valid_point & (angle > 16'd4607 & angle <= 16'd4625);
assign fi_addres[267] = valid_point & (angle > 16'd4625 & angle <= 16'd4634);
assign fi_addres[268] = valid_point & (angle > 16'd4634 & angle <= 16'd4653);
assign fi_addres[269] = valid_point & (angle > 16'd4653 & angle <= 16'd4670);
assign fi_addres[270] = valid_point & (angle > 16'd4670 & angle <= 16'd4688);
assign fi_addres[271] = valid_point & (angle > 16'd4688 & angle <= 16'd4707);
assign fi_addres[272] = valid_point & (angle > 16'd4707 & angle <= 16'd4723);
assign fi_addres[273] = valid_point & (angle > 16'd4723 & angle <= 16'd4741);
assign fi_addres[274] = valid_point & (angle > 16'd4741 & angle <= 16'd4751);
assign fi_addres[275] = valid_point & (angle > 16'd4751 & angle <= 16'd4769);
assign fi_addres[276] = valid_point & (angle > 16'd4769 & angle <= 16'd4787);
assign fi_addres[277] = valid_point & (angle > 16'd4787 & angle <= 16'd4805);
assign fi_addres[278] = valid_point & (angle > 16'd4805 & angle <= 16'd4823);
assign fi_addres[279] = valid_point & (angle > 16'd4823 & angle <= 16'd4841);
assign fi_addres[280] = valid_point & (angle > 16'd4841 & angle <= 16'd4859);
assign fi_addres[281] = valid_point & (angle > 16'd4859 & angle <= 16'd4877);
assign fi_addres[282] = valid_point & (angle > 16'd4877 & angle <= 16'd4886);
assign fi_addres[283] = valid_point & (angle > 16'd4886 & angle <= 16'd4904);
assign fi_addres[284] = valid_point & (angle > 16'd4904 & angle <= 16'd4922);
assign fi_addres[285] = valid_point & (angle > 16'd4922 & angle <= 16'd4940);
assign fi_addres[286] = valid_point & (angle > 16'd4940 & angle <= 16'd4958);
assign fi_addres[287] = valid_point & (angle > 16'd4958 & angle <= 16'd4976);
assign fi_addres[288] = valid_point & (angle > 16'd4976 & angle <= 16'd4994);
assign fi_addres[289] = valid_point & (angle > 16'd4994 & angle <= 16'd5003);
assign fi_addres[290] = valid_point & (angle > 16'd5003 & angle <= 16'd5021);
assign fi_addres[291] = valid_point & (angle > 16'd5021 & angle <= 16'd5039);
assign fi_addres[292] = valid_point & (angle > 16'd5039 & angle <= 16'd5057);
assign fi_addres[293] = valid_point & (angle > 16'd5057 & angle <= 16'd5075);
assign fi_addres[294] = valid_point & (angle > 16'd5075 & angle <= 16'd5093);
assign fi_addres[295] = valid_point & (angle > 16'd5093 & angle <= 16'd5111);
assign fi_addres[296] = valid_point & (angle > 16'd5111 & angle <= 16'd5120);
assign fi_addres[297] = valid_point & (angle > 16'd5120 & angle <= 16'd5138);
assign fi_addres[298] = valid_point & (angle > 16'd5138 & angle <= 16'd5156);
assign fi_addres[299] = valid_point & (angle > 16'd5156 & angle <= 16'd5174);
assign fi_addres[300] = valid_point & (angle > 16'd5174 & angle <= 16'd5192);
assign fi_addres[301] = valid_point & (angle > 16'd5192 & angle <= 16'd5210);
assign fi_addres[302] = valid_point & (angle > 16'd5210 & angle <= 16'd5228);
assign fi_addres[303] = valid_point & (angle > 16'd5228 & angle <= 16'd5237);
assign fi_addres[304] = valid_point & (angle > 16'd5237 & angle <= 16'd5255);
assign fi_addres[305] = valid_point & (angle > 16'd5255 & angle <= 16'd5273);
assign fi_addres[306] = valid_point & (angle > 16'd5273 & angle <= 16'd5291);
assign fi_addres[307] = valid_point & (angle > 16'd5291 & angle <= 16'd5309);
assign fi_addres[308] = valid_point & (angle > 16'd5309 & angle <= 16'd5327);
assign fi_addres[309] = valid_point & (angle > 16'd5327 & angle <= 16'd5345);
assign fi_addres[310] = valid_point & (angle > 16'd5345 & angle <= 16'd5363);
assign fi_addres[311] = valid_point & (angle > 16'd5363 & angle <= 16'd5372);
assign fi_addres[312] = valid_point & (angle > 16'd5372 & angle <= 16'd5390);
assign fi_addres[313] = valid_point & (angle > 16'd5390 & angle <= 16'd5408);
assign fi_addres[314] = valid_point & (angle > 16'd5408 & angle <= 16'd5426);
assign fi_addres[315] = valid_point & (angle > 16'd5426 & angle <= 16'd5444);
assign fi_addres[316] = valid_point & (angle > 16'd5444 & angle <= 16'd5462);
assign fi_addres[317] = valid_point & (angle > 16'd5462 & angle <= 16'd5480);
assign fi_addres[318] = valid_point & (angle > 16'd5480 & angle <= 16'd5489);
assign fi_addres[319] = valid_point & (angle > 16'd5489 & angle <= 16'd5507);
assign fi_addres[320] = valid_point & (angle > 16'd5507 & angle <= 16'd5525);
assign fi_addres[321] = valid_point & (angle > 16'd5525 & angle <= 16'd5543);
assign fi_addres[322] = valid_point & (angle > 16'd5543 & angle <= 16'd5561);
assign fi_addres[323] = valid_point & (angle > 16'd5561 & angle <= 16'd5579);
assign fi_addres[324] = valid_point & (angle > 16'd5579 & angle <= 16'd5597);
assign fi_addres[325] = valid_point & (angle > 16'd5597 & angle <= 16'd5606);
assign fi_addres[326] = valid_point & (angle > 16'd5606 & angle <= 16'd5624);
assign fi_addres[327] = valid_point & (angle > 16'd5624 & angle <= 16'd5642);
assign fi_addres[328] = valid_point & (angle > 16'd5642 & angle <= 16'd5660);
assign fi_addres[329] = valid_point & (angle > 16'd5660 & angle <= 16'd5678);
assign fi_addres[330] = valid_point & (angle > 16'd5678 & angle <= 16'd5696);
assign fi_addres[331] = valid_point & (angle > 16'd5696 & angle <= 16'd5714);
assign fi_addres[332] = valid_point & (angle > 16'd5714 & angle <= 16'd5723);
assign fi_addres[333] = valid_point & (angle > 16'd5723 & angle <= 16'd5741);
assign fi_addres[334] = valid_point & (angle > 16'd5741 & angle <= 16'd5759);
assign fi_addres[335] = valid_point & (angle > 16'd5759 & angle <= 16'd5777);
assign fi_addres[336] = valid_point & (angle > 16'd5777 & angle <= 16'd5795);
assign fi_addres[337] = valid_point & (angle > 16'd5795 & angle <= 16'd5812);
assign fi_addres[338] = valid_point & (angle > 16'd5812 & angle <= 16'd5829);
assign fi_addres[339] = valid_point & (angle > 16'd5829 & angle <= 16'd5848);
assign fi_addres[340] = valid_point & (angle > 16'd5848 & angle <= 16'd5856);
assign fi_addres[341] = valid_point & (angle > 16'd5856 & angle <= 16'd5875);
assign fi_addres[342] = valid_point & (angle > 16'd5875 & angle <= 16'd5892);
assign fi_addres[343] = valid_point & (angle > 16'd5892 & angle <= 16'd5910);
assign fi_addres[344] = valid_point & (angle > 16'd5910 & angle <= 16'd5928);
assign fi_addres[345] = valid_point & (angle > 16'd5928 & angle <= 16'd5946);
assign fi_addres[346] = valid_point & (angle > 16'd5946 & angle <= 16'd5964);
assign fi_addres[347] = valid_point & (angle > 16'd5964 & angle <= 16'd5973);
assign fi_addres[348] = valid_point & (angle > 16'd5973 & angle <= 16'd5991);
assign fi_addres[349] = valid_point & (angle > 16'd5991 & angle <= 16'd6009);
assign fi_addres[350] = valid_point & (angle > 16'd6009 & angle <= 16'd6028);
assign fi_addres[351] = valid_point & (angle > 16'd6028 & angle <= 16'd6045);
assign fi_addres[352] = valid_point & (angle > 16'd6045 & angle <= 16'd6063);
assign fi_addres[353] = valid_point & (angle > 16'd6063 & angle <= 16'd6081);
assign fi_addres[354] = valid_point & (angle > 16'd6081 & angle <= 16'd6090);
assign fi_addres[355] = valid_point & (angle > 16'd6090 & angle <= 16'd6108);
assign fi_addres[356] = valid_point & (angle > 16'd6108 & angle <= 16'd6126);
assign fi_addres[357] = valid_point & (angle > 16'd6126 & angle <= 16'd6144);
assign fi_addres[358] = valid_point & (angle > 16'd6144 & angle <= 16'd6162);
assign fi_addres[359] = valid_point & (angle > 16'd6162 & angle <= 16'd6180);
assign fi_addres[360] = valid_point & (angle > 16'd6180 & angle <= 16'd6198);
assign fi_addres[361] = valid_point & (angle > 16'd6198 & angle <= 16'd6216);
assign fi_addres[362] = valid_point & (angle > 16'd6216 & angle <= 16'd6225);
assign fi_addres[363] = valid_point & (angle > 16'd6225 & angle <= 16'd6243);
assign fi_addres[364] = valid_point & (angle > 16'd6243 & angle <= 16'd6261);
assign fi_addres[365] = valid_point & (angle > 16'd6261 & angle <= 16'd6279);
assign fi_addres[366] = valid_point & (angle > 16'd6279 & angle <= 16'd6297);
assign fi_addres[367] = valid_point & (angle > 16'd6297 & angle <= 16'd6315);
assign fi_addres[368] = valid_point & (angle > 16'd6315 & angle <= 16'd6333);
assign fi_addres[369] = valid_point & (angle > 16'd6333 & angle <= 16'd6342);
assign fi_addres[370] = valid_point & (angle > 16'd6342 & angle <= 16'd6360);
assign fi_addres[371] = valid_point & (angle > 16'd6360 & angle <= 16'd6378);
assign fi_addres[372] = valid_point & (angle > 16'd6378 & angle <= 16'd6396);
assign fi_addres[373] = valid_point & (angle > 16'd6396 & angle <= 16'd6414);
assign fi_addres[374] = valid_point & (angle > 16'd6414 & angle <= 16'd6432);
assign fi_addres[375] = valid_point & (angle > 16'd6432 & angle <= 16'd6450);
assign fi_addres[376] = valid_point & (angle > 16'd6450 & angle <= 16'd6468);
assign fi_addres[377] = valid_point & (angle > 16'd6468 & angle <= 16'd6477);
assign fi_addres[378] = valid_point & (angle > 16'd6477 & angle <= 16'd6495);
assign fi_addres[379] = valid_point & (angle > 16'd6495 & angle <= 16'd6513);
assign fi_addres[380] = valid_point & (angle > 16'd6513 & angle <= 16'd6531);
assign fi_addres[381] = valid_point & (angle > 16'd6531 & angle <= 16'd6549);
assign fi_addres[382] = valid_point & (angle > 16'd6549 & angle <= 16'd6567);
assign fi_addres[383] = valid_point & (angle > 16'd6567 & angle <= 16'd6585);
assign fi_addres[384] = valid_point & (angle > 16'd6585 & angle <= 16'd6594);
assign fi_addres[385] = valid_point & (angle > 16'd6594 & angle <= 16'd6612);
assign fi_addres[386] = valid_point & (angle > 16'd6612 & angle <= 16'd6631);
assign fi_addres[387] = valid_point & (angle > 16'd6631 & angle <= 16'd6648);
assign fi_addres[388] = valid_point & (angle > 16'd6648 & angle <= 16'd6666);
assign fi_addres[389] = valid_point & (angle > 16'd6666 & angle <= 16'd6684);
assign fi_addres[390] = valid_point & (angle > 16'd6684 & angle <= 16'd6702);
assign fi_addres[391] = valid_point & (angle > 16'd6702 & angle <= 16'd6711);
assign fi_addres[392] = valid_point & (angle > 16'd6711 & angle <= 16'd6729);
assign fi_addres[393] = valid_point & (angle > 16'd6729 & angle <= 16'd6747);
assign fi_addres[394] = valid_point & (angle > 16'd6747 & angle <= 16'd6766);
assign fi_addres[395] = valid_point & (angle > 16'd6766 & angle <= 16'd6784);
assign fi_addres[396] = valid_point & (angle > 16'd6784 & angle <= 16'd6802);
assign fi_addres[397] = valid_point & (angle > 16'd6802 & angle <= 16'd6820);
assign fi_addres[398] = valid_point & (angle > 16'd6820 & angle <= 16'd6829);
assign fi_addres[399] = valid_point & (angle > 16'd6829 & angle <= 16'd6847);
assign fi_addres[400] = valid_point & (angle > 16'd6847 & angle <= 16'd6865);
assign fi_addres[401] = valid_point & (angle > 16'd6865 & angle <= 16'd6883);
assign fi_addres[402] = valid_point & (angle > 16'd6883 & angle <= 16'd6901);
assign fi_addres[403] = valid_point & (angle > 16'd6901 & angle <= 16'd6919);
assign fi_addres[404] = valid_point & (angle > 16'd6919 & angle <= 16'd6937);
assign fi_addres[405] = valid_point & (angle > 16'd6937 & angle <= 16'd6955);
assign fi_addres[406] = valid_point & (angle > 16'd6955 & angle <= 16'd6964);
assign fi_addres[407] = valid_point & (angle > 16'd6964 & angle <= 16'd6982);
assign fi_addres[408] = valid_point & (angle > 16'd6982 & angle <= 16'd7000);
assign fi_addres[409] = valid_point & (angle > 16'd7000 & angle <= 16'd7018);
assign fi_addres[410] = valid_point & (angle > 16'd7018 & angle <= 16'd7035);
assign fi_addres[411] = valid_point & (angle > 16'd7035 & angle <= 16'd7052);
assign fi_addres[412] = valid_point & (angle > 16'd7052 & angle <= 16'd7070);
assign fi_addres[413] = valid_point & (angle > 16'd7070 & angle <= 16'd7078);
assign fi_addres[414] = valid_point & (angle > 16'd7078 & angle <= 16'd7096);
assign fi_addres[415] = valid_point & (angle > 16'd7096 & angle <= 16'd7114);
assign fi_addres[416] = valid_point & (angle > 16'd7114 & angle <= 16'd7133);
assign fi_addres[417] = valid_point & (angle > 16'd7133 & angle <= 16'd7151);
assign fi_addres[418] = valid_point & (angle > 16'd7151 & angle <= 16'd7168);
assign fi_addres[419] = valid_point & (angle > 16'd7168 & angle <= 16'd7186);
assign fi_addres[420] = valid_point & (angle > 16'd7186 & angle <= 16'd7196);
assign fi_addres[421] = valid_point & (angle > 16'd7196 & angle <= 16'd7213);
assign fi_addres[422] = valid_point & (angle > 16'd7213 & angle <= 16'd7231);
assign fi_addres[423] = valid_point & (angle > 16'd7231 & angle <= 16'd7250);
assign fi_addres[424] = valid_point & (angle > 16'd7250 & angle <= 16'd7267);
assign fi_addres[425] = valid_point & (angle > 16'd7267 & angle <= 16'd7286);
assign fi_addres[426] = valid_point & (angle > 16'd7286 & angle <= 16'd7304);
assign fi_addres[427] = valid_point & (angle > 16'd7304 & angle <= 16'd7322);
assign fi_addres[428] = valid_point & (angle > 16'd7322 & angle <= 16'd7331);
assign fi_addres[429] = valid_point & (angle > 16'd7331 & angle <= 16'd7351);
assign fi_addres[430] = valid_point & (angle > 16'd7351 & angle <= 16'd7369);
assign fi_addres[431] = valid_point & (angle > 16'd7369 & angle <= 16'd7387);
assign fi_addres[432] = valid_point & (angle > 16'd7387 & angle <= 16'd7405);
assign fi_addres[433] = valid_point & (angle > 16'd7405 & angle <= 16'd7423);
assign fi_addres[434] = valid_point & (angle > 16'd7423 & angle <= 16'd7441);
assign fi_addres[435] = valid_point & (angle > 16'd7441 & angle <= 16'd7450);
assign fi_addres[436] = valid_point & (angle > 16'd7450 & angle <= 16'd7468);
assign fi_addres[437] = valid_point & (angle > 16'd7468 & angle <= 16'd7486);
assign fi_addres[438] = valid_point & (angle > 16'd7486 & angle <= 16'd7504);
assign fi_addres[439] = valid_point & (angle > 16'd7504 & angle <= 16'd7522);
assign fi_addres[440] = valid_point & (angle > 16'd7522 & angle <= 16'd7540);
assign fi_addres[441] = valid_point & (angle > 16'd7540 & angle <= 16'd7558);
assign fi_addres[442] = valid_point & (angle > 16'd7558 & angle <= 16'd7576);
assign fi_addres[443] = valid_point & (angle > 16'd7576 & angle <= 16'd7585);
assign fi_addres[444] = valid_point & (angle > 16'd7585 & angle <= 16'd7603);
assign fi_addres[445] = valid_point & (angle > 16'd7603 & angle <= 16'd7621);
assign fi_addres[446] = valid_point & (angle > 16'd7621 & angle <= 16'd7639);
assign fi_addres[447] = valid_point & (angle > 16'd7639 & angle <= 16'd7657);
assign fi_addres[448] = valid_point & (angle > 16'd7657 & angle <= 16'd7675);
assign fi_addres[449] = valid_point & (angle > 16'd7675 & angle <= 16'd7693);
assign fi_addres[450] = valid_point & (angle > 16'd7693 & angle <= 16'd7702);
assign fi_addres[451] = valid_point & (angle > 16'd7702 & angle <= 16'd7720);
assign fi_addres[452] = valid_point & (angle > 16'd7720 & angle <= 16'd7738);
assign fi_addres[453] = valid_point & (angle > 16'd7738 & angle <= 16'd7756);
assign fi_addres[454] = valid_point & (angle > 16'd7756 & angle <= 16'd7774);
assign fi_addres[455] = valid_point & (angle > 16'd7774 & angle <= 16'd7792);
assign fi_addres[456] = valid_point & (angle > 16'd7792 & angle <= 16'd7810);
assign fi_addres[457] = valid_point & (angle > 16'd7810 & angle <= 16'd7819);
assign fi_addres[458] = valid_point & (angle > 16'd7819 & angle <= 16'd7837);
assign fi_addres[459] = valid_point & (angle > 16'd7837 & angle <= 16'd7853);
assign fi_addres[460] = valid_point & (angle > 16'd7853 & angle <= 16'd7871);
assign fi_addres[461] = valid_point & (angle > 16'd7871 & angle <= 16'd7889);
assign fi_addres[462] = valid_point & (angle > 16'd7889 & angle <= 16'd7907);
assign fi_addres[463] = valid_point & (angle > 16'd7907 & angle <= 16'd7925);
assign fi_addres[464] = valid_point & (angle > 16'd7925 & angle <= 16'd7945);
assign fi_addres[465] = valid_point & (angle > 16'd7945 & angle <= 16'd7954);
assign fi_addres[466] = valid_point & (angle > 16'd7954 & angle <= 16'd7971);
assign fi_addres[467] = valid_point & (angle > 16'd7971 & angle <= 16'd7990);
assign fi_addres[468] = valid_point & (angle > 16'd7990 & angle <= 16'd8008);
assign fi_addres[469] = valid_point & (angle > 16'd8008 & angle <= 16'd8026);
assign fi_addres[470] = valid_point & (angle > 16'd8026 & angle <= 16'd8044);
assign fi_addres[471] = valid_point & (angle > 16'd8044 & angle <= 16'd8062);
assign fi_addres[472] = valid_point & (angle > 16'd8062 & angle <= 16'd8071);
assign fi_addres[473] = valid_point & (angle > 16'd8071 & angle <= 16'd8089);
assign fi_addres[474] = valid_point & (angle > 16'd8089 & angle <= 16'd8107);
assign fi_addres[475] = valid_point & (angle > 16'd8107 & angle <= 16'd8125);
assign fi_addres[476] = valid_point & (angle > 16'd8125 & angle <= 16'd8143);
assign fi_addres[477] = valid_point & (angle > 16'd8143 & angle <= 16'd8161);
assign fi_addres[478] = valid_point & (angle > 16'd8161 & angle <= 16'd8179);
assign fi_addres[479] = valid_point & (angle > 16'd8179 & angle <= 16'd8188);
assign fi_addres[480] = valid_point & (angle > 16'd8188 & angle <= 16'd8206);
assign fi_addres[481] = valid_point & (angle > 16'd8206 & angle <= 16'd8224);
assign fi_addres[482] = valid_point & (angle > 16'd8224 & angle <= 16'd8242);
assign fi_addres[483] = valid_point & (angle > 16'd8242 & angle <= 16'd8260);
assign fi_addres[484] = valid_point & (angle > 16'd8260 & angle <= 16'd8278);
assign fi_addres[485] = valid_point & (angle > 16'd8278 & angle <= 16'd8296);
assign fi_addres[486] = valid_point & (angle > 16'd8296 & angle <= 16'd8314);
assign fi_addres[487] = valid_point & (angle > 16'd8314 & angle <= 16'd8323);
assign fi_addres[488] = valid_point & (angle > 16'd8323 & angle <= 16'd8341);
assign fi_addres[489] = valid_point & (angle > 16'd8341 & angle <= 16'd8359);
assign fi_addres[490] = valid_point & (angle > 16'd8359 & angle <= 16'd8377);
assign fi_addres[491] = valid_point & (angle > 16'd8377 & angle <= 16'd8395);
assign fi_addres[492] = valid_point & (angle > 16'd8395 & angle <= 16'd8413);
assign fi_addres[493] = valid_point & (angle > 16'd8413 & angle <= 16'd8431);
assign fi_addres[494] = valid_point & (angle > 16'd8431 & angle <= 16'd8440);
assign fi_addres[495] = valid_point & (angle > 16'd8440 & angle <= 16'd8458);
assign fi_addres[496] = valid_point & (angle > 16'd8458 & angle <= 16'd8476);
assign fi_addres[497] = valid_point & (angle > 16'd8476 & angle <= 16'd8494);
assign fi_addres[498] = valid_point & (angle > 16'd8494 & angle <= 16'd8512);
assign fi_addres[499] = valid_point & (angle > 16'd8512 & angle <= 16'd8530);
assign fi_addres[500] = valid_point & (angle > 16'd8530 & angle <= 16'd8548);
assign fi_addres[501] = valid_point & (angle > 16'd8548 & angle <= 16'd8557);
assign fi_addres[502] = valid_point & (angle > 16'd8557 & angle <= 16'd8575);
assign fi_addres[503] = valid_point & (angle > 16'd8575 & angle <= 16'd8593);
assign fi_addres[504] = valid_point & (angle > 16'd8593 & angle <= 16'd8611);
assign fi_addres[505] = valid_point & (angle > 16'd8611 & angle <= 16'd8629);
assign fi_addres[506] = valid_point & (angle > 16'd8629 & angle <= 16'd8647);
assign fi_addres[507] = valid_point & (angle > 16'd8647 & angle <= 16'd8665);
assign fi_addres[508] = valid_point & (angle > 16'd8665 & angle <= 16'd8683);
assign fi_addres[509] = valid_point & (angle > 16'd8683 & angle <= 16'd8692);
assign fi_addres[510] = valid_point & (angle > 16'd8692 & angle <= 16'd8710);
assign fi_addres[511] = valid_point & (angle > 16'd8710 & angle <= 16'd8728);
assign fi_addres[512] = valid_point & (angle > 16'd8728 & angle <= 16'd8746);
assign fi_addres[513] = valid_point & (angle > 16'd8746 & angle <= 16'd8764);
assign fi_addres[514] = valid_point & (angle > 16'd8764 & angle <= 16'd8782);
assign fi_addres[515] = valid_point & (angle > 16'd8782 & angle <= 16'd8800);
assign fi_addres[516] = valid_point & (angle > 16'd8800 & angle <= 16'd8809);
assign fi_addres[517] = valid_point & (angle > 16'd8809 & angle <= 16'd8827);
assign fi_addres[518] = valid_point & (angle > 16'd8827 & angle <= 16'd8845);
assign fi_addres[519] = valid_point & (angle > 16'd8845 & angle <= 16'd8863);
assign fi_addres[520] = valid_point & (angle > 16'd8863 & angle <= 16'd8881);
assign fi_addres[521] = valid_point & (angle > 16'd8881 & angle <= 16'd8899);
assign fi_addres[522] = valid_point & (angle > 16'd8899 & angle <= 16'd8917);
assign fi_addres[523] = valid_point & (angle > 16'd8917 & angle <= 16'd8935);
assign fi_addres[524] = valid_point & (angle > 16'd8935 & angle <= 16'd8944);
assign fi_addres[525] = valid_point & (angle > 16'd8944 & angle <= 16'd8962);
assign fi_addres[526] = valid_point & (angle > 16'd8962 & angle <= 16'd8980);
assign fi_addres[527] = valid_point & (angle > 16'd8980 & angle <= 16'd8998);
assign fi_addres[528] = valid_point & (angle > 16'd8998 & angle <= 16'd9016);
assign fi_addres[529] = valid_point & (angle > 16'd9016 & angle <= 16'd9034);
assign fi_addres[530] = valid_point & (angle > 16'd9034 & angle <= 16'd9052);
assign fi_addres[531] = valid_point & (angle > 16'd9052 & angle <= 16'd9061);
assign fi_addres[532] = valid_point & (angle > 16'd9061 & angle <= 16'd9079);
assign fi_addres[533] = valid_point & (angle > 16'd9079 & angle <= 16'd9097);
assign fi_addres[534] = valid_point & (angle > 16'd9097 & angle <= 16'd9115);
assign fi_addres[535] = valid_point & (angle > 16'd9115 & angle <= 16'd9133);
assign fi_addres[536] = valid_point & (angle > 16'd9133 & angle <= 16'd9151);
assign fi_addres[537] = valid_point & (angle > 16'd9151 & angle <= 16'd9169);
assign fi_addres[538] = valid_point & (angle > 16'd9169 & angle <= 16'd9178);
assign fi_addres[539] = valid_point & (angle > 16'd9178 & angle <= 16'd9196);
assign fi_addres[540] = valid_point & (angle > 16'd9196 & angle <= 16'd9214);
assign fi_addres[541] = valid_point & (angle > 16'd9214 & angle <= 16'd9232);
assign fi_addres[542] = valid_point & (angle > 16'd9232 & angle <= 16'd9250);
assign fi_addres[543] = valid_point & (angle > 16'd9250 & angle <= 16'd9268);
assign fi_addres[544] = valid_point & (angle > 16'd9268 & angle <= 16'd9286);
assign fi_addres[545] = valid_point & (angle > 16'd9286 & angle <= 16'd9304);
assign fi_addres[546] = valid_point & (angle > 16'd9304 & angle <= 16'd9315);
assign fi_addres[547] = valid_point & (angle > 16'd9315 & angle <= 16'd9333);
assign fi_addres[548] = valid_point & (angle > 16'd9333 & angle <= 16'd9351);
assign fi_addres[549] = valid_point & (angle > 16'd9351 & angle <= 16'd9369);
assign fi_addres[550] = valid_point & (angle > 16'd9369 & angle <= 16'd9387);
assign fi_addres[551] = valid_point & (angle > 16'd9387 & angle <= 16'd9405);
assign fi_addres[552] = valid_point & (angle > 16'd9405 & angle <= 16'd9423);
assign fi_addres[553] = valid_point & (angle > 16'd9423 & angle <= 16'd9432);
assign fi_addres[554] = valid_point & (angle > 16'd9432 & angle <= 16'd9449);
assign fi_addres[555] = valid_point & (angle > 16'd9449 & angle <= 16'd9467);
assign fi_addres[556] = valid_point & (angle > 16'd9467 & angle <= 16'd9485);
assign fi_addres[557] = valid_point & (angle > 16'd9485 & angle <= 16'd9503);
assign fi_addres[558] = valid_point & (angle > 16'd9503 & angle <= 16'd9521);
assign fi_addres[559] = valid_point & (angle > 16'd9521 & angle <= 16'd9539);
assign fi_addres[560] = valid_point & (angle > 16'd9539 & angle <= 16'd9557);
assign fi_addres[561] = valid_point & (angle > 16'd9557 & angle <= 16'd9566);
assign fi_addres[562] = valid_point & (angle > 16'd9566 & angle <= 16'd9584);
assign fi_addres[563] = valid_point & (angle > 16'd9584 & angle <= 16'd9602);
assign fi_addres[564] = valid_point & (angle > 16'd9602 & angle <= 16'd9619);
assign fi_addres[565] = valid_point & (angle > 16'd9619 & angle <= 16'd9637);
assign fi_addres[566] = valid_point & (angle > 16'd9637 & angle <= 16'd9655);
assign fi_addres[567] = valid_point & (angle > 16'd9655 & angle <= 16'd9673);
assign fi_addres[568] = valid_point & (angle > 16'd9673 & angle <= 16'd9682);
assign fi_addres[569] = valid_point & (angle > 16'd9682 & angle <= 16'd9700);
assign fi_addres[570] = valid_point & (angle > 16'd9700 & angle <= 16'd9718);
assign fi_addres[571] = valid_point & (angle > 16'd9718 & angle <= 16'd9736);
assign fi_addres[572] = valid_point & (angle > 16'd9736 & angle <= 16'd9754);
assign fi_addres[573] = valid_point & (angle > 16'd9754 & angle <= 16'd9772);
assign fi_addres[574] = valid_point & (angle > 16'd9772 & angle <= 16'd9790);
assign fi_addres[575] = valid_point & (angle > 16'd9790 & angle <= 16'd9808);
assign fi_addres[576] = valid_point & (angle > 16'd9808 & angle <= 16'd9817);
assign fi_addres[577] = valid_point & (angle > 16'd9817 & angle <= 16'd9835);
assign fi_addres[578] = valid_point & (angle > 16'd9835 & angle <= 16'd9853);
assign fi_addres[579] = valid_point & (angle > 16'd9853 & angle <= 16'd9871);
assign fi_addres[580] = valid_point & (angle > 16'd9871 & angle <= 16'd9889);
assign fi_addres[581] = valid_point & (angle > 16'd9889 & angle <= 16'd9907);
assign fi_addres[582] = valid_point & (angle > 16'd9907 & angle <= 16'd9925);
assign fi_addres[583] = valid_point & (angle > 16'd9925 & angle <= 16'd9934);
assign fi_addres[584] = valid_point & (angle > 16'd9934 & angle <= 16'd9952);
assign fi_addres[585] = valid_point & (angle > 16'd9952 & angle <= 16'd9970);
assign fi_addres[586] = valid_point & (angle > 16'd9970 & angle <= 16'd9988);
assign fi_addres[587] = valid_point & (angle > 16'd9988 & angle <= 16'd10006);
assign fi_addres[588] = valid_point & (angle > 16'd10006 & angle <= 16'd10024);
assign fi_addres[589] = valid_point & (angle > 16'd10024 & angle <= 16'd10042);
assign fi_addres[590] = valid_point & (angle > 16'd10042 & angle <= 16'd10051);
assign fi_addres[591] = valid_point & (angle > 16'd10051 & angle <= 16'd10069);
assign fi_addres[592] = valid_point & (angle > 16'd10069 & angle <= 16'd10087);
assign fi_addres[593] = valid_point & (angle > 16'd10087 & angle <= 16'd10105);
assign fi_addres[594] = valid_point & (angle > 16'd10105 & angle <= 16'd10123);
assign fi_addres[595] = valid_point & (angle > 16'd10123 & angle <= 16'd10141);
assign fi_addres[596] = valid_point & (angle > 16'd10141 & angle <= 16'd10159);
assign fi_addres[597] = valid_point & (angle > 16'd10159 & angle <= 16'd10177);
assign fi_addres[598] = valid_point & (angle > 16'd10177 & angle <= 16'd10186);
assign fi_addres[599] = valid_point & (angle > 16'd10186 & angle <= 16'd10204);
assign fi_addres[600] = valid_point & (angle > 16'd10204 & angle <= 16'd10222);
assign fi_addres[601] = valid_point & (angle > 16'd10222 & angle <= 16'd10240);
assign fi_addres[602] = valid_point & (angle > 16'd10240 & angle <= 16'd10258);
assign fi_addres[603] = valid_point & (angle > 16'd10258 & angle <= 16'd10276);
assign fi_addres[604] = valid_point & (angle > 16'd10276 & angle <= 16'd10294);
assign fi_addres[605] = valid_point & (angle > 16'd10294 & angle <= 16'd10303);
assign fi_addres[606] = valid_point & (angle > 16'd10303 & angle <= 16'd10321);
assign fi_addres[607] = valid_point & (angle > 16'd10321 & angle <= 16'd10339);
assign fi_addres[608] = valid_point & (angle > 16'd10339 & angle <= 16'd10357);
assign fi_addres[609] = valid_point & (angle > 16'd10357 & angle <= 16'd10375);
assign fi_addres[610] = valid_point & (angle > 16'd10375 & angle <= 16'd10391);
assign fi_addres[611] = valid_point & (angle > 16'd10391 & angle <= 16'd10409);
assign fi_addres[612] = valid_point & (angle > 16'd10409 & angle <= 16'd10418);
assign fi_addres[613] = valid_point & (angle > 16'd10418 & angle <= 16'd10436);
assign fi_addres[614] = valid_point & (angle > 16'd10436 & angle <= 16'd10456);
assign fi_addres[615] = valid_point & (angle > 16'd10456 & angle <= 16'd10474);
assign fi_addres[616] = valid_point & (angle > 16'd10474 & angle <= 16'd10493);
assign fi_addres[617] = valid_point & (angle > 16'd10493 & angle <= 16'd10510);
assign fi_addres[618] = valid_point & (angle > 16'd10510 & angle <= 16'd10528);
assign fi_addres[619] = valid_point & (angle > 16'd10528 & angle <= 16'd10546);
assign fi_addres[620] = valid_point & (angle > 16'd10546 & angle <= 16'd10556);
assign fi_addres[621] = valid_point & (angle > 16'd10556 & angle <= 16'd10574);
assign fi_addres[622] = valid_point & (angle > 16'd10574 & angle <= 16'd10592);
assign fi_addres[623] = valid_point & (angle > 16'd10592 & angle <= 16'd10610);
assign fi_addres[624] = valid_point & (angle > 16'd10610 & angle <= 16'd10628);
assign fi_addres[625] = valid_point & (angle > 16'd10628 & angle <= 16'd10646);
assign fi_addres[626] = valid_point & (angle > 16'd10646 & angle <= 16'd10663);
assign fi_addres[627] = valid_point & (angle > 16'd10663 & angle <= 16'd10672);
assign fi_addres[628] = valid_point & (angle > 16'd10672 & angle <= 16'd10691);
assign fi_addres[629] = valid_point & (angle > 16'd10691 & angle <= 16'd10708);
assign fi_addres[630] = valid_point & (angle > 16'd10708 & angle <= 16'd10726);
assign fi_addres[631] = valid_point & (angle > 16'd10726 & angle <= 16'd10745);
assign fi_addres[632] = valid_point & (angle > 16'd10745 & angle <= 16'd10763);
assign fi_addres[633] = valid_point & (angle > 16'd10763 & angle <= 16'd10781);
assign fi_addres[634] = valid_point & (angle > 16'd10781 & angle <= 16'd10799);
assign fi_addres[635] = valid_point & (angle > 16'd10799 & angle <= 16'd10808);
assign fi_addres[636] = valid_point & (angle > 16'd10808 & angle <= 16'd10826);
assign fi_addres[637] = valid_point & (angle > 16'd10826 & angle <= 16'd10844);
assign fi_addres[638] = valid_point & (angle > 16'd10844 & angle <= 16'd10862);
assign fi_addres[639] = valid_point & (angle > 16'd10862 & angle <= 16'd10880);
assign fi_addres[640] = valid_point & (angle > 16'd10880 & angle <= 16'd10898);
assign fi_addres[641] = valid_point & (angle > 16'd10898 & angle <= 16'd10916);
assign fi_addres[642] = valid_point & (angle > 16'd10916 & angle <= 16'd10925);
assign fi_addres[643] = valid_point & (angle > 16'd10925 & angle <= 16'd10943);
assign fi_addres[644] = valid_point & (angle > 16'd10943 & angle <= 16'd10961);
assign fi_addres[645] = valid_point & (angle > 16'd10961 & angle <= 16'd10979);
assign fi_addres[646] = valid_point & (angle > 16'd10979 & angle <= 16'd10997);
assign fi_addres[647] = valid_point & (angle > 16'd10997 & angle <= 16'd11015);
assign fi_addres[648] = valid_point & (angle > 16'd11015 & angle <= 16'd11033);
assign fi_addres[649] = valid_point & (angle > 16'd11033 & angle <= 16'd11042);
assign fi_addres[650] = valid_point & (angle > 16'd11042 & angle <= 16'd11059);
assign fi_addres[651] = valid_point & (angle > 16'd11059 & angle <= 16'd11077);
assign fi_addres[652] = valid_point & (angle > 16'd11077 & angle <= 16'd11095);
assign fi_addres[653] = valid_point & (angle > 16'd11095 & angle <= 16'd11113);
assign fi_addres[654] = valid_point & (angle > 16'd11113 & angle <= 16'd11132);
assign fi_addres[655] = valid_point & (angle > 16'd11132 & angle <= 16'd11150);
assign fi_addres[656] = valid_point & (angle > 16'd11150 & angle <= 16'd11168);
assign fi_addres[657] = valid_point & (angle > 16'd11168 & angle <= 16'd11177);
assign fi_addres[658] = valid_point & (angle > 16'd11177 & angle <= 16'd11195);
assign fi_addres[659] = valid_point & (angle > 16'd11195 & angle <= 16'd11213);
assign fi_addres[660] = valid_point & (angle > 16'd11213 & angle <= 16'd11231);
assign fi_addres[661] = valid_point & (angle > 16'd11231 & angle <= 16'd11249);
assign fi_addres[662] = valid_point & (angle > 16'd11249 & angle <= 16'd11267);
assign fi_addres[663] = valid_point & (angle > 16'd11267 & angle <= 16'd11285);
assign fi_addres[664] = valid_point & (angle > 16'd11285 & angle <= 16'd11294);
assign fi_addres[665] = valid_point & (angle > 16'd11294 & angle <= 16'd11312);
assign fi_addres[666] = valid_point & (angle > 16'd11312 & angle <= 16'd11330);
assign fi_addres[667] = valid_point & (angle > 16'd11330 & angle <= 16'd11348);
assign fi_addres[668] = valid_point & (angle > 16'd11348 & angle <= 16'd11366);
assign fi_addres[669] = valid_point & (angle > 16'd11366 & angle <= 16'd11384);
assign fi_addres[670] = valid_point & (angle > 16'd11384 & angle <= 16'd11402);
assign fi_addres[671] = valid_point & (angle > 16'd11402 & angle <= 16'd11420);
assign fi_addres[672] = valid_point & (angle > 16'd11420 & angle <= 16'd11429);
assign fi_addres[673] = valid_point & (angle > 16'd11429 & angle <= 16'd11447);
assign fi_addres[674] = valid_point & (angle > 16'd11447 & angle <= 16'd11465);
assign fi_addres[675] = valid_point & (angle > 16'd11465 & angle <= 16'd11483);
assign fi_addres[676] = valid_point & (angle > 16'd11483 & angle <= 16'd11501);
assign fi_addres[677] = valid_point & (angle > 16'd11501 & angle <= 16'd11519);
assign fi_addres[678] = valid_point & (angle > 16'd11519 & angle <= 16'd11537);
assign fi_addres[679] = valid_point & (angle > 16'd11537 & angle <= 16'd11546);
assign fi_addres[680] = valid_point & (angle > 16'd11546 & angle <= 16'd11564);
assign fi_addres[681] = valid_point & (angle > 16'd11564 & angle <= 16'd11582);
assign fi_addres[682] = valid_point & (angle > 16'd11582 & angle <= 16'd11600);
assign fi_addres[683] = valid_point & (angle > 16'd11600 & angle <= 16'd11618);
assign fi_addres[684] = valid_point & (angle > 16'd11618 & angle <= 16'd11637);
assign fi_addres[685] = valid_point & (angle > 16'd11637 & angle <= 16'd11655);
assign fi_addres[686] = valid_point & (angle > 16'd11655 & angle <= 16'd11672);
assign fi_addres[687] = valid_point & (angle > 16'd11672 & angle <= 16'd11681);
assign fi_addres[688] = valid_point & (angle > 16'd11681 & angle <= 16'd11700);
assign fi_addres[689] = valid_point & (angle > 16'd11700 & angle <= 16'd11718);
assign fi_addres[690] = valid_point & (angle > 16'd11718 & angle <= 16'd11735);
assign fi_addres[691] = valid_point & (angle > 16'd11735 & angle <= 16'd11753);
assign fi_addres[692] = valid_point & (angle > 16'd11753 & angle <= 16'd11771);
assign fi_addres[693] = valid_point & (angle > 16'd11771 & angle <= 16'd11789);
assign fi_addres[694] = valid_point & (angle > 16'd11789 & angle <= 16'd11798);
assign fi_addres[695] = valid_point & (angle > 16'd11798 & angle <= 16'd11816);
assign fi_addres[696] = valid_point & (angle > 16'd11816 & angle <= 16'd11835);
assign fi_addres[697] = valid_point & (angle > 16'd11835 & angle <= 16'd11852);
assign fi_addres[698] = valid_point & (angle > 16'd11852 & angle <= 16'd11870);
assign fi_addres[699] = valid_point & (angle > 16'd11870 & angle <= 16'd11888);
assign fi_addres[700] = valid_point & (angle > 16'd11888 & angle <= 16'd11906);
assign fi_addres[701] = valid_point & (angle > 16'd11906 & angle <= 16'd11924);
assign fi_addres[702] = valid_point & (angle > 16'd11924 & angle <= 16'd11933);
assign fi_addres[703] = valid_point & (angle > 16'd11933 & angle <= 16'd11951);
assign fi_addres[704] = valid_point & (angle > 16'd11951 & angle <= 16'd11969);
assign fi_addres[705] = valid_point & (angle > 16'd11969 & angle <= 16'd11987);
assign fi_addres[706] = valid_point & (angle > 16'd11987 & angle <= 16'd12005);
assign fi_addres[707] = valid_point & (angle > 16'd12005 & angle <= 16'd12023);
assign fi_addres[708] = valid_point & (angle > 16'd12023 & angle <= 16'd12041);
assign fi_addres[709] = valid_point & (angle > 16'd12041 & angle <= 16'd12050);
assign fi_addres[710] = valid_point & (angle > 16'd12050 & angle <= 16'd12068);
assign fi_addres[711] = valid_point & (angle > 16'd12068 & angle <= 16'd12086);
assign fi_addres[712] = valid_point & (angle > 16'd12086 & angle <= 16'd12104);
assign fi_addres[713] = valid_point & (angle > 16'd12104 & angle <= 16'd12122);
assign fi_addres[714] = valid_point & (angle > 16'd12122 & angle <= 16'd12140);
assign fi_addres[715] = valid_point & (angle > 16'd12140 & angle <= 16'd12158);
assign fi_addres[716] = valid_point & (angle > 16'd12158 & angle <= 16'd12176);
assign fi_addres[717] = valid_point & (angle > 16'd12176 & angle <= 16'd12185);
assign fi_addres[718] = valid_point & (angle > 16'd12185 & angle <= 16'd12203);
assign fi_addres[719] = valid_point & (angle > 16'd12203 & angle <= 16'd12221);
assign fi_addres[720] = valid_point & (angle > 16'd12221 & angle <= 16'd12239);
assign fi_addres[721] = valid_point & (angle > 16'd12239 & angle <= 16'd12257);
assign fi_addres[722] = valid_point & (angle > 16'd12257 & angle <= 16'd12275);
assign fi_addres[723] = valid_point & (angle > 16'd12275 & angle <= 16'd12293);
assign fi_addres[724] = valid_point & (angle > 16'd12293 & angle <= 16'd12302);
assign fi_addres[725] = valid_point & (angle > 16'd12302 & angle <= 16'd12320);
assign fi_addres[726] = valid_point & (angle > 16'd12320 & angle <= 16'd12338);
assign fi_addres[727] = valid_point & (angle > 16'd12338 & angle <= 16'd12356);
assign fi_addres[728] = valid_point & (angle > 16'd12356 & angle <= 16'd12374);
assign fi_addres[729] = valid_point & (angle > 16'd12374 & angle <= 16'd12392);
assign fi_addres[730] = valid_point & (angle > 16'd12392 & angle <= 16'd12410);
assign fi_addres[731] = valid_point & (angle > 16'd12410 & angle <= 16'd12419);
assign fi_addres[732] = valid_point & (angle > 16'd12419 & angle <= 16'd12437);
assign fi_addres[733] = valid_point & (angle > 16'd12437 & angle <= 16'd12455);
assign fi_addres[734] = valid_point & (angle > 16'd12455 & angle <= 16'd12473);
assign fi_addres[735] = valid_point & (angle > 16'd12473 & angle <= 16'd12491);
assign fi_addres[736] = valid_point & (angle > 16'd12491 & angle <= 16'd12509);
assign fi_addres[737] = valid_point & (angle > 16'd12509 & angle <= 16'd12527);
assign fi_addres[738] = valid_point & (angle > 16'd12527 & angle <= 16'd12545);
assign fi_addres[739] = valid_point & (angle > 16'd12545 & angle <= 16'd12554);
assign fi_addres[740] = valid_point & (angle > 16'd12554 & angle <= 16'd12572);
assign fi_addres[741] = valid_point & (angle > 16'd12572 & angle <= 16'd12590);
assign fi_addres[742] = valid_point & (angle > 16'd12590 & angle <= 16'd12608);
assign fi_addres[743] = valid_point & (angle > 16'd12608 & angle <= 16'd12626);
assign fi_addres[744] = valid_point & (angle > 16'd12626 & angle <= 16'd12644);
assign fi_addres[745] = valid_point & (angle > 16'd12644 & angle <= 16'd12662);
assign fi_addres[746] = valid_point & (angle > 16'd12662 & angle <= 16'd12680);
assign fi_addres[747] = valid_point & (angle > 16'd12680 & angle <= 16'd12689);
assign fi_addres[748] = valid_point & (angle > 16'd12689 & angle <= 16'd12708);
assign fi_addres[749] = valid_point & (angle > 16'd12708 & angle <= 16'd12726);
assign fi_addres[750] = valid_point & (angle > 16'd12726 & angle <= 16'd12743);
assign fi_addres[751] = valid_point & (angle > 16'd12743 & angle <= 16'd12762);
assign fi_addres[752] = valid_point & (angle > 16'd12762 & angle <= 16'd12780);
assign fi_addres[753] = valid_point & (angle > 16'd12780 & angle <= 16'd12797);
assign fi_addres[754] = valid_point & (angle > 16'd12797 & angle <= 16'd12807);
assign fi_addres[755] = valid_point & (angle > 16'd12807 & angle <= 16'd12825);
assign fi_addres[756] = valid_point & (angle > 16'd12825 & angle <= 16'd12843);
assign fi_addres[757] = valid_point & (angle > 16'd12843 & angle <= 16'd12861);
assign fi_addres[758] = valid_point & (angle > 16'd12861 & angle <= 16'd12879);
assign fi_addres[759] = valid_point & (angle > 16'd12879 & angle <= 16'd12897);
assign fi_addres[760] = valid_point & (angle > 16'd12897 & angle <= 16'd12915);
assign fi_addres[761] = valid_point & (angle > 16'd12915 & angle <= 16'd12922);
assign fi_addres[762] = valid_point & (angle > 16'd12922 & angle <= 16'd12940);
assign fi_addres[763] = valid_point & (angle > 16'd12940 & angle <= 16'd12958);
assign fi_addres[764] = valid_point & (angle > 16'd12958 & angle <= 16'd12976);
assign fi_addres[765] = valid_point & (angle > 16'd12976 & angle <= 16'd12994);
assign fi_addres[766] = valid_point & (angle > 16'd12994 & angle <= 16'd13012);
assign fi_addres[767] = valid_point & (angle > 16'd13012 & angle <= 16'd13030);
assign fi_addres[768] = valid_point & (angle > 16'd13030 & angle <= 16'd13048);
assign fi_addres[769] = valid_point & (angle > 16'd13048 & angle <= 16'd13059);
assign fi_addres[770] = valid_point & (angle > 16'd13059 & angle <= 16'd13077);
assign fi_addres[771] = valid_point & (angle > 16'd13077 & angle <= 16'd13095);
assign fi_addres[772] = valid_point & (angle > 16'd13095 & angle <= 16'd13113);
assign fi_addres[773] = valid_point & (angle > 16'd13113 & angle <= 16'd13131);
assign fi_addres[774] = valid_point & (angle > 16'd13131 & angle <= 16'd13149);
assign fi_addres[775] = valid_point & (angle > 16'd13149 & angle <= 16'd13167);
assign fi_addres[776] = valid_point & (angle > 16'd13167 & angle <= 16'd13176);
assign fi_addres[777] = valid_point & (angle > 16'd13176 & angle <= 16'd13194);
assign fi_addres[778] = valid_point & (angle > 16'd13194 & angle <= 16'd13212);
assign fi_addres[779] = valid_point & (angle > 16'd13212 & angle <= 16'd13230);
assign fi_addres[780] = valid_point & (angle > 16'd13230 & angle <= 16'd13248);
assign fi_addres[781] = valid_point & (angle > 16'd13248 & angle <= 16'd13266);
assign fi_addres[782] = valid_point & (angle > 16'd13266 & angle <= 16'd13287);
assign fi_addres[783] = valid_point & (angle > 16'd13287 & angle <= 16'd13305);
assign fi_addres[784] = valid_point & (angle > 16'd13305 & angle <= 16'd13314);
assign fi_addres[785] = valid_point & (angle > 16'd13314 & angle <= 16'd13332);
assign fi_addres[786] = valid_point & (angle > 16'd13332 & angle <= 16'd13350);
assign fi_addres[787] = valid_point & (angle > 16'd13350 & angle <= 16'd13368);
assign fi_addres[788] = valid_point & (angle > 16'd13368 & angle <= 16'd13386);
assign fi_addres[789] = valid_point & (angle > 16'd13386 & angle <= 16'd13404);
assign fi_addres[790] = valid_point & (angle > 16'd13404 & angle <= 16'd13422);
assign fi_addres[791] = valid_point & (angle > 16'd13422 & angle <= 16'd13431);
assign fi_addres[792] = valid_point & (angle > 16'd13431 & angle <= 16'd13449);
assign fi_addres[793] = valid_point & (angle > 16'd13449 & angle <= 16'd13467);
assign fi_addres[794] = valid_point & (angle > 16'd13467 & angle <= 16'd13485);
assign fi_addres[795] = valid_point & (angle > 16'd13485 & angle <= 16'd13503);
assign fi_addres[796] = valid_point & (angle > 16'd13503 & angle <= 16'd13521);
assign fi_addres[797] = valid_point & (angle > 16'd13521 & angle <= 16'd13539);
assign fi_addres[798] = valid_point & (angle > 16'd13539 & angle <= 16'd13557);
assign fi_addres[799] = valid_point & (angle > 16'd13557 & angle <= 16'd13566);
assign fi_addres[800] = valid_point & (angle > 16'd13566 & angle <= 16'd13584);
assign fi_addres[801] = valid_point & (angle > 16'd13584 & angle <= 16'd13602);
assign fi_addres[802] = valid_point & (angle > 16'd13602 & angle <= 16'd13620);
assign fi_addres[803] = valid_point & (angle > 16'd13620 & angle <= 16'd13638);
assign fi_addres[804] = valid_point & (angle > 16'd13638 & angle <= 16'd13656);
assign fi_addres[805] = valid_point & (angle > 16'd13656 & angle <= 16'd13674);
assign fi_addres[806] = valid_point & (angle > 16'd13674 & angle <= 16'd13682);
assign fi_addres[807] = valid_point & (angle > 16'd13682 & angle <= 16'd13701);
assign fi_addres[808] = valid_point & (angle > 16'd13701 & angle <= 16'd13718);
assign fi_addres[809] = valid_point & (angle > 16'd13718 & angle <= 16'd13736);
assign fi_addres[810] = valid_point & (angle > 16'd13736 & angle <= 16'd13754);
assign fi_addres[811] = valid_point & (angle > 16'd13754 & angle <= 16'd13772);
assign fi_addres[812] = valid_point & (angle > 16'd13772 & angle <= 16'd13790);
assign fi_addres[813] = valid_point & (angle > 16'd13790 & angle <= 16'd13799);
assign fi_addres[814] = valid_point & (angle > 16'd13799 & angle <= 16'd13817);
assign fi_addres[815] = valid_point & (angle > 16'd13817 & angle <= 16'd13835);
assign fi_addres[816] = valid_point & (angle > 16'd13835 & angle <= 16'd13853);
assign fi_addres[817] = valid_point & (angle > 16'd13853 & angle <= 16'd13871);
assign fi_addres[818] = valid_point & (angle > 16'd13871 & angle <= 16'd13889);
assign fi_addres[819] = valid_point & (angle > 16'd13889 & angle <= 16'd13907);
assign fi_addres[820] = valid_point & (angle > 16'd13907 & angle <= 16'd13925);
assign fi_addres[821] = valid_point & (angle > 16'd13925 & angle <= 16'd13953);
assign fi_addres[822] = valid_point & (angle > 16'd13953 & angle <= 16'd13971);
assign fi_addres[823] = valid_point & (angle > 16'd13971 & angle <= 16'd14003);
assign fi_addres[824] = valid_point & (angle > 16'd14003 & angle <= 16'd14021);
assign fi_addres[825] = valid_point & (angle > 16'd14021 & angle <= 16'd14039);
assign fi_addres[826] = valid_point & (angle > 16'd14039 & angle <= 16'd14052);
assign fi_addres[827] = valid_point & (angle > 16'd14052 & angle <= 16'd14084);
assign fi_addres[828] = valid_point & (angle > 16'd14084 & angle <= 16'd14102);
assign fi_addres[829] = valid_point & (angle > 16'd14102 & angle <= 16'd14121);
assign fi_addres[830] = valid_point & (angle > 16'd14121 & angle <= 16'd14141);
assign fi_addres[831] = valid_point & (angle > 16'd14141 & angle <= 16'd14159);
assign fi_addres[832] = valid_point & (angle > 16'd14159 & angle <= 16'd14177);
assign fi_addres[833] = valid_point & (angle > 16'd14177 & angle <= 16'd14186);
assign fi_addres[834] = valid_point & (angle > 16'd14186 & angle <= 16'd14204);
assign fi_addres[835] = valid_point & (angle > 16'd14204 & angle <= 16'd14222);
assign fi_addres[836] = valid_point & (angle > 16'd14222 & angle <= 16'd14241);
assign fi_addres[837] = valid_point & (angle > 16'd14241 & angle <= 16'd14259);
assign fi_addres[838] = valid_point & (angle > 16'd14259 & angle <= 16'd14276);
assign fi_addres[839] = valid_point & (angle > 16'd14276 & angle <= 16'd14295);
assign fi_addres[840] = valid_point & (angle > 16'd14295 & angle <= 16'd14304);
assign fi_addres[841] = valid_point & (angle > 16'd14304 & angle <= 16'd14322);
assign fi_addres[842] = valid_point & (angle > 16'd14322 & angle <= 16'd14340);
assign fi_addres[843] = valid_point & (angle > 16'd14340 & angle <= 16'd14358);
assign fi_addres[844] = valid_point & (angle > 16'd14358 & angle <= 16'd14375);
assign fi_addres[845] = valid_point & (angle > 16'd14375 & angle <= 16'd14394);
assign fi_addres[846] = valid_point & (angle > 16'd14394 & angle <= 16'd14411);
assign fi_addres[847] = valid_point & (angle > 16'd14411 & angle <= 16'd14421);
assign fi_addres[848] = valid_point & (angle > 16'd14421 & angle <= 16'd14438);
assign fi_addres[849] = valid_point & (angle > 16'd14438 & angle <= 16'd14456);
assign fi_addres[850] = valid_point & (angle > 16'd14456 & angle <= 16'd14474);
assign fi_addres[851] = valid_point & (angle > 16'd14474 & angle <= 16'd14492);
assign fi_addres[852] = valid_point & (angle > 16'd14492 & angle <= 16'd14510);
assign fi_addres[853] = valid_point & (angle > 16'd14510 & angle <= 16'd14528);
assign fi_addres[854] = valid_point & (angle > 16'd14528 & angle <= 16'd14546);
assign fi_addres[855] = valid_point & (angle > 16'd14546 & angle <= 16'd14555);
assign fi_addres[856] = valid_point & (angle > 16'd14555 & angle <= 16'd14574);
assign fi_addres[857] = valid_point & (angle > 16'd14574 & angle <= 16'd14591);
assign fi_addres[858] = valid_point & (angle > 16'd14591 & angle <= 16'd14609);
assign fi_addres[859] = valid_point & (angle > 16'd14609 & angle <= 16'd14627);
assign fi_addres[860] = valid_point & (angle > 16'd14627 & angle <= 16'd14645);
assign fi_addres[861] = valid_point & (angle > 16'd14645 & angle <= 16'd14664);
assign fi_addres[862] = valid_point & (angle > 16'd14664 & angle <= 16'd14672);
assign fi_addres[863] = valid_point & (angle > 16'd14672 & angle <= 16'd14690);
assign fi_addres[864] = valid_point & (angle > 16'd14690 & angle <= 16'd14708);
assign fi_addres[865] = valid_point & (angle > 16'd14708 & angle <= 16'd14726);
assign fi_addres[866] = valid_point & (angle > 16'd14726 & angle <= 16'd14745);
assign fi_addres[867] = valid_point & (angle > 16'd14745 & angle <= 16'd14762);
assign fi_addres[868] = valid_point & (angle > 16'd14762 & angle <= 16'd14780);
assign fi_addres[869] = valid_point & (angle > 16'd14780 & angle <= 16'd14790);
assign fi_addres[870] = valid_point & (angle > 16'd14790 & angle <= 16'd14808);
assign fi_addres[871] = valid_point & (angle > 16'd14808 & angle <= 16'd14825);
assign fi_addres[872] = valid_point & (angle > 16'd14825 & angle <= 16'd14844);
assign fi_addres[873] = valid_point & (angle > 16'd14844 & angle <= 16'd14862);
assign fi_addres[874] = valid_point & (angle > 16'd14862 & angle <= 16'd14880);
assign fi_addres[875] = valid_point & (angle > 16'd14880 & angle <= 16'd14897);
assign fi_addres[876] = valid_point & (angle > 16'd14897 & angle <= 16'd14916);
assign fi_addres[877] = valid_point & (angle > 16'd14916 & angle <= 16'd14924);
assign fi_addres[878] = valid_point & (angle > 16'd14924 & angle <= 16'd14943);
assign fi_addres[879] = valid_point & (angle > 16'd14943 & angle <= 16'd14960);
assign fi_addres[880] = valid_point & (angle > 16'd14960 & angle <= 16'd14978);
assign fi_addres[881] = valid_point & (angle > 16'd14978 & angle <= 16'd14996);
assign fi_addres[882] = valid_point & (angle > 16'd14996 & angle <= 16'd15014);
assign fi_addres[883] = valid_point & (angle > 16'd15014 & angle <= 16'd15032);
assign fi_addres[884] = valid_point & (angle > 16'd15032 & angle <= 16'd15041);
assign fi_addres[885] = valid_point & (angle > 16'd15041 & angle <= 16'd15059);
assign fi_addres[886] = valid_point & (angle > 16'd15059 & angle <= 16'd15077);
assign fi_addres[887] = valid_point & (angle > 16'd15077 & angle <= 16'd15096);
assign fi_addres[888] = valid_point & (angle > 16'd15096 & angle <= 16'd15114);
assign fi_addres[889] = valid_point & (angle > 16'd15114 & angle <= 16'd15131);
assign fi_addres[890] = valid_point & (angle > 16'd15131 & angle <= 16'd15149);
assign fi_addres[891] = valid_point & (angle > 16'd15149 & angle <= 16'd15167);
assign fi_addres[892] = valid_point & (angle > 16'd15167 & angle <= 16'd15176);
assign fi_addres[893] = valid_point & (angle > 16'd15176 & angle <= 16'd15194);
assign fi_addres[894] = valid_point & (angle > 16'd15194 & angle <= 16'd15212);
assign fi_addres[895] = valid_point & (angle > 16'd15212 & angle <= 16'd15230);
assign fi_addres[896] = valid_point & (angle > 16'd15230 & angle <= 16'd15248);
assign fi_addres[897] = valid_point & (angle > 16'd15248 & angle <= 16'd15267);
assign fi_addres[898] = valid_point & (angle > 16'd15267 & angle <= 16'd15284);
assign fi_addres[899] = valid_point & (angle > 16'd15284 & angle <= 16'd15294);
assign fi_addres[900] = valid_point & (angle > 16'd15294 & angle <= 16'd15311);
assign fi_addres[901] = valid_point & (angle > 16'd15311 & angle <= 16'd15329);
assign fi_addres[902] = valid_point & (angle > 16'd15329 & angle <= 16'd15347);
assign fi_addres[903] = valid_point & (angle > 16'd15347 & angle <= 16'd15365);
assign fi_addres[904] = valid_point & (angle > 16'd15365 & angle <= 16'd15383);
assign fi_addres[905] = valid_point & (angle > 16'd15383 & angle <= 16'd15401);
assign fi_addres[906] = valid_point & (angle > 16'd15401 & angle <= 16'd15410);
assign fi_addres[907] = valid_point & (angle > 16'd15410 & angle <= 16'd15429);
assign fi_addres[908] = valid_point & (angle > 16'd15429 & angle <= 16'd15447);
assign fi_addres[909] = valid_point & (angle > 16'd15447 & angle <= 16'd15464);
assign fi_addres[910] = valid_point & (angle > 16'd15464 & angle <= 16'd15483);
assign fi_addres[911] = valid_point & (angle > 16'd15483 & angle <= 16'd15501);
assign fi_addres[912] = valid_point & (angle > 16'd15501 & angle <= 16'd15519);
assign fi_addres[913] = valid_point & (angle > 16'd15519 & angle <= 16'd15528);
assign fi_addres[914] = valid_point & (angle > 16'd15528 & angle <= 16'd15546);
assign fi_addres[915] = valid_point & (angle > 16'd15546 & angle <= 16'd15564);
assign fi_addres[916] = valid_point & (angle > 16'd15564 & angle <= 16'd15582);
assign fi_addres[917] = valid_point & (angle > 16'd15582 & angle <= 16'd15600);
assign fi_addres[918] = valid_point & (angle > 16'd15600 & angle <= 16'd15617);
assign fi_addres[919] = valid_point & (angle > 16'd15617 & angle <= 16'd15635);
assign fi_addres[920] = valid_point & (angle > 16'd15635 & angle <= 16'd15653);
assign fi_addres[921] = valid_point & (angle > 16'd15653 & angle <= 16'd15662);
assign fi_addres[922] = valid_point & (angle > 16'd15662 & angle <= 16'd15680);
assign fi_addres[923] = valid_point & (angle > 16'd15680 & angle <= 16'd15698);
assign fi_addres[924] = valid_point & (angle > 16'd15698 & angle <= 16'd15716);
assign fi_addres[925] = valid_point & (angle > 16'd15716 & angle <= 16'd15734);
assign fi_addres[926] = valid_point & (angle > 16'd15734 & angle <= 16'd15752);
assign fi_addres[927] = valid_point & (angle > 16'd15752 & angle <= 16'd15770);
assign fi_addres[928] = valid_point & (angle > 16'd15770 & angle <= 16'd15789);
assign fi_addres[929] = valid_point & (angle > 16'd15789 & angle <= 16'd15797);
assign fi_addres[930] = valid_point & (angle > 16'd15797 & angle <= 16'd15816);
assign fi_addres[931] = valid_point & (angle > 16'd15816 & angle <= 16'd15834);
assign fi_addres[932] = valid_point & (angle > 16'd15834 & angle <= 16'd15852);
assign fi_addres[933] = valid_point & (angle > 16'd15852 & angle <= 16'd15869);
assign fi_addres[934] = valid_point & (angle > 16'd15869 & angle <= 16'd15888);
assign fi_addres[935] = valid_point & (angle > 16'd15888 & angle <= 16'd15906);
assign fi_addres[936] = valid_point & (angle > 16'd15906 & angle <= 16'd15914);
assign fi_addres[937] = valid_point & (angle > 16'd15914 & angle <= 16'd15932);
assign fi_addres[938] = valid_point & (angle > 16'd15932 & angle <= 16'd15950);
assign fi_addres[939] = valid_point & (angle > 16'd15950 & angle <= 16'd15969);
assign fi_addres[940] = valid_point & (angle > 16'd15969 & angle <= 16'd15987);
assign fi_addres[941] = valid_point & (angle > 16'd15987 & angle <= 16'd16005);
assign fi_addres[942] = valid_point & (angle > 16'd16005 & angle <= 16'd16023);
assign fi_addres[943] = valid_point & (angle > 16'd16023 & angle <= 16'd16032);
assign fi_addres[944] = valid_point & (angle > 16'd16032 & angle <= 16'd16049);
assign fi_addres[945] = valid_point & (angle > 16'd16049 & angle <= 16'd16067);
assign fi_addres[946] = valid_point & (angle > 16'd16067 & angle <= 16'd16085);
assign fi_addres[947] = valid_point & (angle > 16'd16085 & angle <= 16'd16104);
assign fi_addres[948] = valid_point & (angle > 16'd16104 & angle <= 16'd16122);
assign fi_addres[949] = valid_point & (angle > 16'd16122 & angle <= 16'd16140);
assign fi_addres[950] = valid_point & (angle > 16'd16140 & angle <= 16'd16149);
assign fi_addres[951] = valid_point & (angle > 16'd16149 & angle <= 16'd16167);
assign fi_addres[952] = valid_point & (angle > 16'd16167 & angle <= 16'd16185);
assign fi_addres[953] = valid_point & (angle > 16'd16185 & angle <= 16'd16203);
assign fi_addres[954] = valid_point & (angle > 16'd16203 & angle <= 16'd16221);
assign fi_addres[955] = valid_point & (angle > 16'd16221 & angle <= 16'd16239);
assign fi_addres[956] = valid_point & (angle > 16'd16239 & angle <= 16'd16266);
assign fi_addres[957] = valid_point & (angle > 16'd16266 & angle <= 16'd16296);
assign fi_addres[958] = valid_point & (angle > 16'd16296 & angle <= 16'd16324);
assign fi_addres[959] = valid_point & (angle > 16'd16324 & angle <= 16'd16342);
assign fi_addres[960] = valid_point & (angle > 16'd16342 & angle <= 16'd16360);
assign fi_addres[961] = valid_point & (angle > 16'd16360 & angle <= 16'd16378);
assign fi_addres[962] = valid_point & (angle > 16'd16378 & angle <= 16'd16396);
assign fi_addres[963] = valid_point & (angle > 16'd16396 & angle <= 16'd16413);
assign fi_addres[964] = valid_point & (angle > 16'd16413 & angle <= 16'd16430);
assign fi_addres[965] = valid_point & (angle > 16'd16430 & angle <= 16'd16448);
assign fi_addres[966] = valid_point & (angle > 16'd16448 & angle <= 16'd16471);
assign fi_addres[967] = valid_point & (angle > 16'd16471 & angle <= 16'd16491);
assign fi_addres[968] = valid_point & (angle > 16'd16491 & angle <= 16'd16509);
assign fi_addres[969] = valid_point & (angle > 16'd16509 & angle <= 16'd16518);
assign fi_addres[970] = valid_point & (angle > 16'd16518 & angle <= 16'd16536);
assign fi_addres[971] = valid_point & (angle > 16'd16536 & angle <= 16'd16554);
assign fi_addres[972] = valid_point & (angle > 16'd16554 & angle <= 16'd16572);
assign fi_addres[973] = valid_point & (angle > 16'd16572 & angle <= 16'd16590);
assign fi_addres[974] = valid_point & (angle > 16'd16590 & angle <= 16'd16608);
assign fi_addres[975] = valid_point & (angle > 16'd16608 & angle <= 16'd16626);
assign fi_addres[976] = valid_point & (angle > 16'd16626 & angle <= 16'd16635);
assign fi_addres[977] = valid_point & (angle > 16'd16635 & angle <= 16'd16653);
assign fi_addres[978] = valid_point & (angle > 16'd16653 & angle <= 16'd16671);
assign fi_addres[979] = valid_point & (angle > 16'd16671 & angle <= 16'd16689);
assign fi_addres[980] = valid_point & (angle > 16'd16689 & angle <= 16'd16708);
assign fi_addres[981] = valid_point & (angle > 16'd16708 & angle <= 16'd16727);
assign fi_addres[982] = valid_point & (angle > 16'd16727 & angle <= 16'd16756);
assign fi_addres[983] = valid_point & (angle > 16'd16756 & angle <= 16'd16774);
assign fi_addres[984] = valid_point & (angle > 16'd16774 & angle <= 16'd16792);
assign fi_addres[985] = valid_point & (angle > 16'd16792 & angle <= 16'd16822);
assign fi_addres[986] = valid_point & (angle > 16'd16822 & angle <= 16'd16840);
assign fi_addres[987] = valid_point & (angle > 16'd16840 & angle <= 16'd16857);
assign fi_addres[988] = valid_point & (angle > 16'd16857 & angle <= 16'd16884);
assign fi_addres[989] = valid_point & (angle > 16'd16884 & angle <= 16'd16902);
assign fi_addres[990] = valid_point & (angle > 16'd16902 & angle <= 16'd16920);
assign fi_addres[991] = valid_point & (angle > 16'd16920 & angle <= 16'd16938);
assign fi_addres[992] = valid_point & (angle > 16'd16938 & angle <= 16'd16955);
assign fi_addres[993] = valid_point & (angle > 16'd16955 & angle <= 16'd16972);
assign fi_addres[994] = valid_point & (angle > 16'd16972 & angle <= 16'd16990);
assign fi_addres[995] = valid_point & (angle > 16'd16990 & angle <= 16'd17017);
assign fi_addres[996] = valid_point & (angle > 16'd17017 & angle <= 16'd17035);
assign fi_addres[997] = valid_point & (angle > 16'd17035 & angle <= 16'd17053);
assign fi_addres[998] = valid_point & (angle > 16'd17053 & angle <= 16'd17079);
assign fi_addres[999] = valid_point & (angle > 16'd17079 & angle <= 16'd17097);
assign fi_addres[1000] = valid_point & (angle > 16'd17097 & angle <= 16'd17118);
assign fi_addres[1001] = valid_point & (angle > 16'd17118 & angle <= 16'd17136);
assign fi_addres[1002] = valid_point & (angle > 16'd17136 & angle <= 16'd17154);
assign fi_addres[1003] = valid_point & (angle > 16'd17154 & angle <= 16'd17172);
assign fi_addres[1004] = valid_point & (angle > 16'd17172 & angle <= 16'd17190);
assign fi_addres[1005] = valid_point & (angle > 16'd17190 & angle <= 16'd17208);
assign fi_addres[1006] = valid_point & (angle > 16'd17208 & angle <= 16'd17236);
assign fi_addres[1007] = valid_point & (angle > 16'd17236 & angle <= 16'd17253);
assign fi_addres[1008] = valid_point & (angle > 16'd17253 & angle <= 16'd17271);
assign fi_addres[1009] = valid_point & (angle > 16'd17271 & angle <= 16'd17289);
assign fi_addres[1010] = valid_point & (angle > 16'd17289 & angle <= 16'd17307);
assign fi_addres[1011] = valid_point & (angle > 16'd17307 & angle <= 16'd17325);
assign fi_addres[1012] = valid_point & (angle > 16'd17325 & angle <= 16'd17349);
assign fi_addres[1013] = valid_point & (angle > 16'd17349 & angle <= 16'd17367);
assign fi_addres[1014] = valid_point & (angle > 16'd17367 & angle <= 16'd17395);
assign fi_addres[1015] = valid_point & (angle > 16'd17395 & angle <= 16'd17424);
assign fi_addres[1016] = valid_point & (angle > 16'd17424 & angle <= 16'd17442);
assign fi_addres[1017] = valid_point & (angle > 16'd17442 & angle <= 16'd17460);
assign fi_addres[1018] = valid_point & (angle > 16'd17460 & angle <= 16'd17478);
assign fi_addres[1019] = valid_point & (angle > 16'd17478 & angle <= 16'd17505);
assign fi_addres[1020] = valid_point & (angle > 16'd17505 & angle <= 16'd17523);
assign fi_addres[1021] = valid_point & (angle > 16'd17523 & angle <= 16'd17541);
assign fi_addres[1022] = valid_point & (angle > 16'd17541 & angle <= 16'd17559);
assign fi_addres[1023] = valid_point & (angle > 16'd17559 & angle <= 16'd17577);
assign fi_addres[1024] = valid_point & (angle > 16'd17577 & angle <= 16'd17595);
assign fi_addres[1025] = valid_point & (angle > 16'd17595 & angle <= 16'd17613);
assign fi_addres[1026] = valid_point & (angle > 16'd17613 & angle <= 16'd17640);
assign fi_addres[1027] = valid_point & (angle > 16'd17640 & angle <= 16'd17658);
assign fi_addres[1028] = valid_point & (angle > 16'd17658 & angle <= 16'd17676);
assign fi_addres[1029] = valid_point & (angle > 16'd17676 & angle <= 16'd17694);
assign fi_addres[1030] = valid_point & (angle > 16'd17694 & angle <= 16'd17719);
assign fi_addres[1031] = valid_point & (angle > 16'd17719 & angle <= 16'd17737);
assign fi_addres[1032] = valid_point & (angle > 16'd17737 & angle <= 16'd17764);
assign fi_addres[1033] = valid_point & (angle > 16'd17764 & angle <= 16'd17793);
assign fi_addres[1034] = valid_point & (angle > 16'd17793 & angle <= 16'd17821);
assign fi_addres[1035] = valid_point & (angle > 16'd17821 & angle <= 16'd17847);
assign fi_addres[1036] = valid_point & (angle > 16'd17847 & angle <= 16'd17874);
assign fi_addres[1037] = valid_point & (angle > 16'd17874 & angle <= 16'd17900);
assign fi_addres[1038] = valid_point & (angle > 16'd17900 & angle <= 16'd17917);
assign fi_addres[1039] = valid_point & (angle > 16'd17917 & angle <= 16'd17935);
assign fi_addres[1040] = valid_point & (angle > 16'd17935 & angle <= 16'd17964);
assign fi_addres[1041] = valid_point & (angle > 16'd17964 & angle <= 16'd17982);
assign fi_addres[1042] = valid_point & (angle > 16'd17982 & angle <= 16'd18009);
assign fi_addres[1043] = valid_point & (angle > 16'd18009 & angle <= 16'd18035);
assign fi_addres[1044] = valid_point & (angle > 16'd18035 & angle <= 16'd18063);
assign fi_addres[1045] = valid_point & (angle > 16'd18063 & angle <= 16'd18089);
assign fi_addres[1046] = valid_point & (angle > 16'd18089 & angle <= 16'd18108);
assign fi_addres[1047] = valid_point & (angle > 16'd18108 & angle <= 16'd18126);
assign fi_addres[1048] = valid_point & (angle > 16'd18126 & angle <= 16'd18154);
assign fi_addres[1049] = valid_point & (angle > 16'd18154 & angle <= 16'd18180);
assign fi_addres[1050] = valid_point & (angle > 16'd18180 & angle <= 16'd18198);
assign fi_addres[1051] = valid_point & (angle > 16'd18198 & angle <= 16'd18224);
assign fi_addres[1052] = valid_point & (angle > 16'd18224 & angle <= 16'd18251);
assign fi_addres[1053] = valid_point & (angle > 16'd18251 & angle <= 16'd18269);
assign fi_addres[1054] = valid_point & (angle > 16'd18269 & angle <= 16'd18287);
assign fi_addres[1055] = valid_point & (angle > 16'd18287 & angle <= 16'd18315);
assign fi_addres[1056] = valid_point & (angle > 16'd18315 & angle <= 16'd18333);
assign fi_addres[1057] = valid_point & (angle > 16'd18333 & angle <= 16'd18351);
assign fi_addres[1058] = valid_point & (angle > 16'd18351 & angle <= 16'd18368);
assign fi_addres[1059] = valid_point & (angle > 16'd18368 & angle <= 16'd18386);
assign fi_addres[1060] = valid_point & (angle > 16'd18386 & angle <= 16'd18403);
assign fi_addres[1061] = valid_point & (angle > 16'd18403 & angle <= 16'd18422);
assign fi_addres[1062] = valid_point & (angle > 16'd18422 & angle <= 16'd18442);
assign fi_addres[1063] = valid_point & (angle > 16'd18442 & angle <= 16'd18469);
assign fi_addres[1064] = valid_point & (angle > 16'd18469 & angle <= 16'd18487);
assign fi_addres[1065] = valid_point & (angle > 16'd18487 & angle <= 16'd18504);
assign fi_addres[1066] = valid_point & (angle > 16'd18504 & angle <= 16'd18523);
assign fi_addres[1067] = valid_point & (angle > 16'd18523 & angle <= 16'd18541);
assign fi_addres[1068] = valid_point & (angle > 16'd18541 & angle <= 16'd18558);
assign fi_addres[1069] = valid_point & (angle > 16'd18558 & angle <= 16'd18575);
assign fi_addres[1070] = valid_point & (angle > 16'd18575 & angle <= 16'd18592);
assign fi_addres[1071] = valid_point & (angle > 16'd18592 & angle <= 16'd18621);
assign fi_addres[1072] = valid_point & (angle > 16'd18621 & angle <= 16'd18640);
assign fi_addres[1073] = valid_point & (angle > 16'd18640 & angle <= 16'd18658);
assign fi_addres[1074] = valid_point & (angle > 16'd18658 & angle <= 16'd18691);
assign fi_addres[1075] = valid_point & (angle > 16'd18691 & angle <= 16'd18710);
assign fi_addres[1076] = valid_point & (angle > 16'd18710 & angle <= 16'd18737);
assign fi_addres[1077] = valid_point & (angle > 16'd18737 & angle <= 16'd18756);
assign fi_addres[1078] = valid_point & (angle > 16'd18756 & angle <= 16'd18775);
assign fi_addres[1079] = valid_point & (angle > 16'd18775 & angle <= 16'd18793);
assign fi_addres[1080] = valid_point & (angle > 16'd18793 & angle <= 16'd18811);
assign fi_addres[1081] = valid_point & (angle > 16'd18811 & angle <= 16'd18838);
assign fi_addres[1082] = valid_point & (angle > 16'd18838 & angle <= 16'd18856);
assign fi_addres[1083] = valid_point & (angle > 16'd18856 & angle <= 16'd18874);
assign fi_addres[1084] = valid_point & (angle > 16'd18874 & angle <= 16'd18891);
assign fi_addres[1085] = valid_point & (angle > 16'd18891 & angle <= 16'd18917);
assign fi_addres[1086] = valid_point & (angle > 16'd18917 & angle <= 16'd18935);
assign fi_addres[1087] = valid_point & (angle > 16'd18935 & angle <= 16'd18953);
assign fi_addres[1088] = valid_point & (angle > 16'd18953 & angle <= 16'd18971);
assign fi_addres[1089] = valid_point & (angle > 16'd18971 & angle <= 16'd18989);
assign fi_addres[1090] = valid_point & (angle > 16'd18989 & angle <= 16'd19016);
assign fi_addres[1091] = valid_point & (angle > 16'd19016 & angle <= 16'd19047);
assign fi_addres[1092] = valid_point & (angle > 16'd19047 & angle <= 16'd19068);
assign fi_addres[1093] = valid_point & (angle > 16'd19068 & angle <= 16'd19096);
assign fi_addres[1094] = valid_point & (angle > 16'd19096 & angle <= 16'd19114);
assign fi_addres[1095] = valid_point & (angle > 16'd19114 & angle <= 16'd19133);
assign fi_addres[1096] = valid_point & (angle > 16'd19133 & angle <= 16'd19151);
assign fi_addres[1097] = valid_point & (angle > 16'd19151 & angle <= 16'd19169);
assign fi_addres[1098] = valid_point & (angle > 16'd19169 & angle <= 16'd19187);
assign fi_addres[1099] = valid_point & (angle > 16'd19187 & angle <= 16'd19207);
assign fi_addres[1100] = valid_point & (angle > 16'd19207 & angle <= 16'd19223);
assign fi_addres[1101] = valid_point & (angle > 16'd19223 & angle <= 16'd19241);
assign fi_addres[1102] = valid_point & (angle > 16'd19241 & angle <= 16'd19257);
assign fi_addres[1103] = valid_point & (angle > 16'd19257 & angle <= 16'd19274);
assign fi_addres[1104] = valid_point & (angle > 16'd19274 & angle <= 16'd19299);
assign fi_addres[1105] = valid_point & (angle > 16'd19299 & angle <= 16'd19317);
assign fi_addres[1106] = valid_point & (angle > 16'd19317 & angle <= 16'd19335);
assign fi_addres[1107] = valid_point & (angle > 16'd19335 & angle <= 16'd19353);
assign fi_addres[1108] = valid_point & (angle > 16'd19353 & angle <= 16'd19362);
assign fi_addres[1109] = valid_point & (angle > 16'd19362 & angle <= 16'd19380);
assign fi_addres[1110] = valid_point & (angle > 16'd19380 & angle <= 16'd19398);
assign fi_addres[1111] = valid_point & (angle > 16'd19398 & angle <= 16'd19416);
assign fi_addres[1112] = valid_point & (angle > 16'd19416 & angle <= 16'd19434);
assign fi_addres[1113] = valid_point & (angle > 16'd19434 & angle <= 16'd19452);
assign fi_addres[1114] = valid_point & (angle > 16'd19452 & angle <= 16'd19470);
assign fi_addres[1115] = valid_point & (angle > 16'd19470 & angle <= 16'd19488);
assign fi_addres[1116] = valid_point & (angle > 16'd19488 & angle <= 16'd19497);
assign fi_addres[1117] = valid_point & (angle > 16'd19497 & angle <= 16'd19515);
assign fi_addres[1118] = valid_point & (angle > 16'd19515 & angle <= 16'd19533);
assign fi_addres[1119] = valid_point & (angle > 16'd19533 & angle <= 16'd19551);
assign fi_addres[1120] = valid_point & (angle > 16'd19551 & angle <= 16'd19569);
assign fi_addres[1121] = valid_point & (angle > 16'd19569 & angle <= 16'd19587);
assign fi_addres[1122] = valid_point & (angle > 16'd19587 & angle <= 16'd19605);
assign fi_addres[1123] = valid_point & (angle > 16'd19605 & angle <= 16'd19615);
assign fi_addres[1124] = valid_point & (angle > 16'd19615 & angle <= 16'd19632);
assign fi_addres[1125] = valid_point & (angle > 16'd19632 & angle <= 16'd19650);
assign fi_addres[1126] = valid_point & (angle > 16'd19650 & angle <= 16'd19668);
assign fi_addres[1127] = valid_point & (angle > 16'd19668 & angle <= 16'd19686);
assign fi_addres[1128] = valid_point & (angle > 16'd19686 & angle <= 16'd19704);
assign fi_addres[1129] = valid_point & (angle > 16'd19704 & angle <= 16'd19728);
assign fi_addres[1130] = valid_point & (angle > 16'd19728 & angle <= 16'd19749);
assign fi_addres[1131] = valid_point & (angle > 16'd19749 & angle <= 16'd19767);
assign fi_addres[1132] = valid_point & (angle > 16'd19767 & angle <= 16'd19785);
assign fi_addres[1133] = valid_point & (angle > 16'd19785 & angle <= 16'd19803);
assign fi_addres[1134] = valid_point & (angle > 16'd19803 & angle <= 16'd19821);
assign fi_addres[1135] = valid_point & (angle > 16'd19821 & angle <= 16'd19839);
assign fi_addres[1136] = valid_point & (angle > 16'd19839 & angle <= 16'd19848);
assign fi_addres[1137] = valid_point & (angle > 16'd19848 & angle <= 16'd19866);
assign fi_addres[1138] = valid_point & (angle > 16'd19866 & angle <= 16'd19884);
assign fi_addres[1139] = valid_point & (angle > 16'd19884 & angle <= 16'd19902);
assign fi_addres[1140] = valid_point & (angle > 16'd19902 & angle <= 16'd19920);
assign fi_addres[1141] = valid_point & (angle > 16'd19920 & angle <= 16'd19938);
assign fi_addres[1142] = valid_point & (angle > 16'd19938 & angle <= 16'd19956);
assign fi_addres[1143] = valid_point & (angle > 16'd19956 & angle <= 16'd19974);
assign fi_addres[1144] = valid_point & (angle > 16'd19974 & angle <= 16'd19983);
assign fi_addres[1145] = valid_point & (angle > 16'd19983 & angle <= 16'd20001);
assign fi_addres[1146] = valid_point & (angle > 16'd20001 & angle <= 16'd20019);
assign fi_addres[1147] = valid_point & (angle > 16'd20019 & angle <= 16'd20037);
assign fi_addres[1148] = valid_point & (angle > 16'd20037 & angle <= 16'd20055);
assign fi_addres[1149] = valid_point & (angle > 16'd20055 & angle <= 16'd20073);
assign fi_addres[1150] = valid_point & (angle > 16'd20073 & angle <= 16'd20091);
assign fi_addres[1151] = valid_point & (angle > 16'd20091 & angle <= 16'd20100);
assign fi_addres[1152] = valid_point & (angle > 16'd20100 & angle <= 16'd20118);
assign fi_addres[1153] = valid_point & (angle > 16'd20118 & angle <= 16'd20136);
assign fi_addres[1154] = valid_point & (angle > 16'd20136 & angle <= 16'd20154);
assign fi_addres[1155] = valid_point & (angle > 16'd20154 & angle <= 16'd20172);
assign fi_addres[1156] = valid_point & (angle > 16'd20172 & angle <= 16'd20190);
assign fi_addres[1157] = valid_point & (angle > 16'd20190 & angle <= 16'd20208);
assign fi_addres[1158] = valid_point & (angle > 16'd20208 & angle <= 16'd20226);
assign fi_addres[1159] = valid_point & (angle > 16'd20226 & angle <= 16'd20235);
assign fi_addres[1160] = valid_point & (angle > 16'd20235 & angle <= 16'd20253);
assign fi_addres[1161] = valid_point & (angle > 16'd20253 & angle <= 16'd20271);
assign fi_addres[1162] = valid_point & (angle > 16'd20271 & angle <= 16'd20289);
assign fi_addres[1163] = valid_point & (angle > 16'd20289 & angle <= 16'd20307);
assign fi_addres[1164] = valid_point & (angle > 16'd20307 & angle <= 16'd20325);
assign fi_addres[1165] = valid_point & (angle > 16'd20325 & angle <= 16'd20343);
assign fi_addres[1166] = valid_point & (angle > 16'd20343 & angle <= 16'd20352);
assign fi_addres[1167] = valid_point & (angle > 16'd20352 & angle <= 16'd20370);
assign fi_addres[1168] = valid_point & (angle > 16'd20370 & angle <= 16'd20388);
assign fi_addres[1169] = valid_point & (angle > 16'd20388 & angle <= 16'd20406);
assign fi_addres[1170] = valid_point & (angle > 16'd20406 & angle <= 16'd20424);
assign fi_addres[1171] = valid_point & (angle > 16'd20424 & angle <= 16'd20442);
assign fi_addres[1172] = valid_point & (angle > 16'd20442 & angle <= 16'd20460);
assign fi_addres[1173] = valid_point & (angle > 16'd20460 & angle <= 16'd20469);
assign fi_addres[1174] = valid_point & (angle > 16'd20469 & angle <= 16'd20487);
assign fi_addres[1175] = valid_point & (angle > 16'd20487 & angle <= 16'd20504);
assign fi_addres[1176] = valid_point & (angle > 16'd20504 & angle <= 16'd20522);
assign fi_addres[1177] = valid_point & (angle > 16'd20522 & angle <= 16'd20540);
assign fi_addres[1178] = valid_point & (angle > 16'd20540 & angle <= 16'd20558);
assign fi_addres[1179] = valid_point & (angle > 16'd20558 & angle <= 16'd20576);
assign fi_addres[1180] = valid_point & (angle > 16'd20576 & angle <= 16'd20585);
assign fi_addres[1181] = valid_point & (angle > 16'd20585 & angle <= 16'd20603);
assign fi_addres[1182] = valid_point & (angle > 16'd20603 & angle <= 16'd20621);
assign fi_addres[1183] = valid_point & (angle > 16'd20621 & angle <= 16'd20639);
assign fi_addres[1184] = valid_point & (angle > 16'd20639 & angle <= 16'd20657);
assign fi_addres[1185] = valid_point & (angle > 16'd20657 & angle <= 16'd20675);
assign fi_addres[1186] = valid_point & (angle > 16'd20675 & angle <= 16'd20693);
assign fi_addres[1187] = valid_point & (angle > 16'd20693 & angle <= 16'd20711);
assign fi_addres[1188] = valid_point & (angle > 16'd20711 & angle <= 16'd20734);
assign fi_addres[1189] = valid_point & (angle > 16'd20734 & angle <= 16'd20755);
assign fi_addres[1190] = valid_point & (angle > 16'd20755 & angle <= 16'd20773);
assign fi_addres[1191] = valid_point & (angle > 16'd20773 & angle <= 16'd20791);
assign fi_addres[1192] = valid_point & (angle > 16'd20791 & angle <= 16'd20809);
assign fi_addres[1193] = valid_point & (angle > 16'd20809 & angle <= 16'd20827);
assign fi_addres[1194] = valid_point & (angle > 16'd20827 & angle <= 16'd20836);
assign fi_addres[1195] = valid_point & (angle > 16'd20836 & angle <= 16'd20854);
assign fi_addres[1196] = valid_point & (angle > 16'd20854 & angle <= 16'd20872);
assign fi_addres[1197] = valid_point & (angle > 16'd20872 & angle <= 16'd20890);
assign fi_addres[1198] = valid_point & (angle > 16'd20890 & angle <= 16'd20907);
assign fi_addres[1199] = valid_point & (angle > 16'd20907 & angle <= 16'd20925);
assign fi_addres[1200] = valid_point & (angle > 16'd20925 & angle <= 16'd20943);
assign fi_addres[1201] = valid_point & (angle > 16'd20943 & angle <= 16'd20961);
assign fi_addres[1202] = valid_point & (angle > 16'd20961 & angle <= 16'd20970);
assign fi_addres[1203] = valid_point & (angle > 16'd20970 & angle <= 16'd20988);
assign fi_addres[1204] = valid_point & (angle > 16'd20988 & angle <= 16'd21006);
assign fi_addres[1205] = valid_point & (angle > 16'd21006 & angle <= 16'd21024);
assign fi_addres[1206] = valid_point & (angle > 16'd21024 & angle <= 16'd21042);
assign fi_addres[1207] = valid_point & (angle > 16'd21042 & angle <= 16'd21060);
assign fi_addres[1208] = valid_point & (angle > 16'd21060 & angle <= 16'd21078);
assign fi_addres[1209] = valid_point & (angle > 16'd21078 & angle <= 16'd21087);
assign fi_addres[1210] = valid_point & (angle > 16'd21087 & angle <= 16'd21105);
assign fi_addres[1211] = valid_point & (angle > 16'd21105 & angle <= 16'd21123);
assign fi_addres[1212] = valid_point & (angle > 16'd21123 & angle <= 16'd21141);
assign fi_addres[1213] = valid_point & (angle > 16'd21141 & angle <= 16'd21159);
assign fi_addres[1214] = valid_point & (angle > 16'd21159 & angle <= 16'd21177);
assign fi_addres[1215] = valid_point & (angle > 16'd21177 & angle <= 16'd21195);
assign fi_addres[1216] = valid_point & (angle > 16'd21195 & angle <= 16'd21204);
assign fi_addres[1217] = valid_point & (angle > 16'd21204 & angle <= 16'd21222);
assign fi_addres[1218] = valid_point & (angle > 16'd21222 & angle <= 16'd21240);
assign fi_addres[1219] = valid_point & (angle > 16'd21240 & angle <= 16'd21258);
assign fi_addres[1220] = valid_point & (angle > 16'd21258 & angle <= 16'd21276);
assign fi_addres[1221] = valid_point & (angle > 16'd21276 & angle <= 16'd21294);
assign fi_addres[1222] = valid_point & (angle > 16'd21294 & angle <= 16'd21312);
assign fi_addres[1223] = valid_point & (angle > 16'd21312 & angle <= 16'd21330);
assign fi_addres[1224] = valid_point & (angle > 16'd21330 & angle <= 16'd21339);
assign fi_addres[1225] = valid_point & (angle > 16'd21339 & angle <= 16'd21357);
assign fi_addres[1226] = valid_point & (angle > 16'd21357 & angle <= 16'd21375);
assign fi_addres[1227] = valid_point & (angle > 16'd21375 & angle <= 16'd21393);
assign fi_addres[1228] = valid_point & (angle > 16'd21393 & angle <= 16'd21411);
assign fi_addres[1229] = valid_point & (angle > 16'd21411 & angle <= 16'd21429);
assign fi_addres[1230] = valid_point & (angle > 16'd21429 & angle <= 16'd21447);
assign fi_addres[1231] = valid_point & (angle > 16'd21447 & angle <= 16'd21455);
assign fi_addres[1232] = valid_point & (angle > 16'd21455 & angle <= 16'd21473);
assign fi_addres[1233] = valid_point & (angle > 16'd21473 & angle <= 16'd21492);
assign fi_addres[1234] = valid_point & (angle > 16'd21492 & angle <= 16'd21509);
assign fi_addres[1235] = valid_point & (angle > 16'd21509 & angle <= 16'd21527);
assign fi_addres[1236] = valid_point & (angle > 16'd21527 & angle <= 16'd21545);
assign fi_addres[1237] = valid_point & (angle > 16'd21545 & angle <= 16'd21563);
assign fi_addres[1238] = valid_point & (angle > 16'd21563 & angle <= 16'd21572);
assign fi_addres[1239] = valid_point & (angle > 16'd21572 & angle <= 16'd21590);
assign fi_addres[1240] = valid_point & (angle > 16'd21590 & angle <= 16'd21608);
assign fi_addres[1241] = valid_point & (angle > 16'd21608 & angle <= 16'd21626);
assign fi_addres[1242] = valid_point & (angle > 16'd21626 & angle <= 16'd21644);
assign fi_addres[1243] = valid_point & (angle > 16'd21644 & angle <= 16'd21662);
assign fi_addres[1244] = valid_point & (angle > 16'd21662 & angle <= 16'd21680);
assign fi_addres[1245] = valid_point & (angle > 16'd21680 & angle <= 16'd21689);
assign fi_addres[1246] = valid_point & (angle > 16'd21689 & angle <= 16'd21707);
assign fi_addres[1247] = valid_point & (angle > 16'd21707 & angle <= 16'd21725);
assign fi_addres[1248] = valid_point & (angle > 16'd21725 & angle <= 16'd21743);
assign fi_addres[1249] = valid_point & (angle > 16'd21743 & angle <= 16'd21761);
assign fi_addres[1250] = valid_point & (angle > 16'd21761 & angle <= 16'd21779);
assign fi_addres[1251] = valid_point & (angle > 16'd21779 & angle <= 16'd21797);
assign fi_addres[1252] = valid_point & (angle > 16'd21797 & angle <= 16'd21806);
assign fi_addres[1253] = valid_point & (angle > 16'd21806 & angle <= 16'd21824);
assign fi_addres[1254] = valid_point & (angle > 16'd21824 & angle <= 16'd21842);
assign fi_addres[1255] = valid_point & (angle > 16'd21842 & angle <= 16'd21860);
assign fi_addres[1256] = valid_point & (angle > 16'd21860 & angle <= 16'd21878);
assign fi_addres[1257] = valid_point & (angle > 16'd21878 & angle <= 16'd21896);
assign fi_addres[1258] = valid_point & (angle > 16'd21896 & angle <= 16'd21914);
assign fi_addres[1259] = valid_point & (angle > 16'd21914 & angle <= 16'd21932);
assign fi_addres[1260] = valid_point & (angle > 16'd21932 & angle <= 16'd21941);
assign fi_addres[1261] = valid_point & (angle > 16'd21941 & angle <= 16'd21959);
assign fi_addres[1262] = valid_point & (angle > 16'd21959 & angle <= 16'd21977);
assign fi_addres[1263] = valid_point & (angle > 16'd21977 & angle <= 16'd21995);
assign fi_addres[1264] = valid_point & (angle > 16'd21995 & angle <= 16'd22013);
assign fi_addres[1265] = valid_point & (angle > 16'd22013 & angle <= 16'd22031);
assign fi_addres[1266] = valid_point & (angle > 16'd22031 & angle <= 16'd22048);
assign fi_addres[1267] = valid_point & (angle > 16'd22048 & angle <= 16'd22057);
assign fi_addres[1268] = valid_point & (angle > 16'd22057 & angle <= 16'd22075);
assign fi_addres[1269] = valid_point & (angle > 16'd22075 & angle <= 16'd22094);
assign fi_addres[1270] = valid_point & (angle > 16'd22094 & angle <= 16'd22111);
assign fi_addres[1271] = valid_point & (angle > 16'd22111 & angle <= 16'd22129);
assign fi_addres[1272] = valid_point & (angle > 16'd22129 & angle <= 16'd22147);
assign fi_addres[1273] = valid_point & (angle > 16'd22147 & angle <= 16'd22165);
assign fi_addres[1274] = valid_point & (angle > 16'd22165 & angle <= 16'd22174);
assign fi_addres[1275] = valid_point & (angle > 16'd22174 & angle <= 16'd22192);
assign fi_addres[1276] = valid_point & (angle > 16'd22192 & angle <= 16'd22210);
assign fi_addres[1277] = valid_point & (angle > 16'd22210 & angle <= 16'd22228);
assign fi_addres[1278] = valid_point & (angle > 16'd22228 & angle <= 16'd22246);
assign fi_addres[1279] = valid_point & (angle > 16'd22246 & angle <= 16'd22264);
assign fi_addres[1280] = valid_point & (angle > 16'd22264 & angle <= 16'd22282);
assign fi_addres[1281] = valid_point & (angle > 16'd22282 & angle <= 16'd22300);
assign fi_addres[1282] = valid_point & (angle > 16'd22300 & angle <= 16'd22309);
assign fi_addres[1283] = valid_point & (angle > 16'd22309 & angle <= 16'd22327);
assign fi_addres[1284] = valid_point & (angle > 16'd22327 & angle <= 16'd22345);
assign fi_addres[1285] = valid_point & (angle > 16'd22345 & angle <= 16'd22363);
assign fi_addres[1286] = valid_point & (angle > 16'd22363 & angle <= 16'd22381);
assign fi_addres[1287] = valid_point & (angle > 16'd22381 & angle <= 16'd22399);
assign fi_addres[1288] = valid_point & (angle > 16'd22399 & angle <= 16'd22417);
assign fi_addres[1289] = valid_point & (angle > 16'd22417 & angle <= 16'd22426);
assign fi_addres[1290] = valid_point & (angle > 16'd22426 & angle <= 16'd22444);
assign fi_addres[1291] = valid_point & (angle > 16'd22444 & angle <= 16'd22462);
assign fi_addres[1292] = valid_point & (angle > 16'd22462 & angle <= 16'd22480);
assign fi_addres[1293] = valid_point & (angle > 16'd22480 & angle <= 16'd22498);
assign fi_addres[1294] = valid_point & (angle > 16'd22498 & angle <= 16'd22516);
assign fi_addres[1295] = valid_point & (angle > 16'd22516 & angle <= 16'd22534);
assign fi_addres[1296] = valid_point & (angle > 16'd22534 & angle <= 16'd22552);
assign fi_addres[1297] = valid_point & (angle > 16'd22552 & angle <= 16'd22561);
assign fi_addres[1298] = valid_point & (angle > 16'd22561 & angle <= 16'd22579);
assign fi_addres[1299] = valid_point & (angle > 16'd22579 & angle <= 16'd22597);
assign fi_addres[1300] = valid_point & (angle > 16'd22597 & angle <= 16'd22615);
assign fi_addres[1301] = valid_point & (angle > 16'd22615 & angle <= 16'd22633);
assign fi_addres[1302] = valid_point & (angle > 16'd22633 & angle <= 16'd22651);
assign fi_addres[1303] = valid_point & (angle > 16'd22651 & angle <= 16'd22669);
assign fi_addres[1304] = valid_point & (angle > 16'd22669 & angle <= 16'd22678);
assign fi_addres[1305] = valid_point & (angle > 16'd22678 & angle <= 16'd22696);
assign fi_addres[1306] = valid_point & (angle > 16'd22696 & angle <= 16'd22714);
assign fi_addres[1307] = valid_point & (angle > 16'd22714 & angle <= 16'd22732);
assign fi_addres[1308] = valid_point & (angle > 16'd22732 & angle <= 16'd22750);
assign fi_addres[1309] = valid_point & (angle > 16'd22750 & angle <= 16'd22768);
assign fi_addres[1310] = valid_point & (angle > 16'd22768 & angle <= 16'd22786);
assign fi_addres[1311] = valid_point & (angle > 16'd22786 & angle <= 16'd22795);
assign fi_addres[1312] = valid_point & (angle > 16'd22795 & angle <= 16'd22813);
assign fi_addres[1313] = valid_point & (angle > 16'd22813 & angle <= 16'd22831);
assign fi_addres[1314] = valid_point & (angle > 16'd22831 & angle <= 16'd22849);
assign fi_addres[1315] = valid_point & (angle > 16'd22849 & angle <= 16'd22867);
assign fi_addres[1316] = valid_point & (angle > 16'd22867 & angle <= 16'd22885);
assign fi_addres[1317] = valid_point & (angle > 16'd22885 & angle <= 16'd22902);
assign fi_addres[1318] = valid_point & (angle > 16'd22902 & angle <= 16'd22911);
assign fi_addres[1319] = valid_point & (angle > 16'd22911 & angle <= 16'd22930);
assign fi_addres[1320] = valid_point & (angle > 16'd22930 & angle <= 16'd22948);
assign fi_addres[1321] = valid_point & (angle > 16'd22948 & angle <= 16'd22966);
assign fi_addres[1322] = valid_point & (angle > 16'd22966 & angle <= 16'd22984);
assign fi_addres[1323] = valid_point & (angle > 16'd22984 & angle <= 16'd23002);
assign fi_addres[1324] = valid_point & (angle > 16'd23002 & angle <= 16'd23019);
assign fi_addres[1325] = valid_point & (angle > 16'd23019 & angle <= 16'd23028);
assign fi_addres[1326] = valid_point & (angle > 16'd23028 & angle <= 16'd23047);
assign fi_addres[1327] = valid_point & (angle > 16'd23047 & angle <= 16'd23064);
assign fi_addres[1328] = valid_point & (angle > 16'd23064 & angle <= 16'd23083);
assign fi_addres[1329] = valid_point & (angle > 16'd23083 & angle <= 16'd23100);
assign fi_addres[1330] = valid_point & (angle > 16'd23100 & angle <= 16'd23118);
assign fi_addres[1331] = valid_point & (angle > 16'd23118 & angle <= 16'd23136);
assign fi_addres[1332] = valid_point & (angle > 16'd23136 & angle <= 16'd23154);
assign fi_addres[1333] = valid_point & (angle > 16'd23154 & angle <= 16'd23163);
assign fi_addres[1334] = valid_point & (angle > 16'd23163 & angle <= 16'd23181);
assign fi_addres[1335] = valid_point & (angle > 16'd23181 & angle <= 16'd23199);
assign fi_addres[1336] = valid_point & (angle > 16'd23199 & angle <= 16'd23217);
assign fi_addres[1337] = valid_point & (angle > 16'd23217 & angle <= 16'd23235);
assign fi_addres[1338] = valid_point & (angle > 16'd23235 & angle <= 16'd23253);
assign fi_addres[1339] = valid_point & (angle > 16'd23253 & angle <= 16'd23271);
assign fi_addres[1340] = valid_point & (angle > 16'd23271 & angle <= 16'd23280);
assign fi_addres[1341] = valid_point & (angle > 16'd23280 & angle <= 16'd23298);
assign fi_addres[1342] = valid_point & (angle > 16'd23298 & angle <= 16'd23316);
assign fi_addres[1343] = valid_point & (angle > 16'd23316 & angle <= 16'd23334);
assign fi_addres[1344] = valid_point & (angle > 16'd23334 & angle <= 16'd23352);
assign fi_addres[1345] = valid_point & (angle > 16'd23352 & angle <= 16'd23370);
assign fi_addres[1346] = valid_point & (angle > 16'd23370 & angle <= 16'd23388);
assign fi_addres[1347] = valid_point & (angle > 16'd23388 & angle <= 16'd23397);
assign fi_addres[1348] = valid_point & (angle > 16'd23397 & angle <= 16'd23415);
assign fi_addres[1349] = valid_point & (angle > 16'd23415 & angle <= 16'd23433);
assign fi_addres[1350] = valid_point & (angle > 16'd23433 & angle <= 16'd23451);
assign fi_addres[1351] = valid_point & (angle > 16'd23451 & angle <= 16'd23469);
assign fi_addres[1352] = valid_point & (angle > 16'd23469 & angle <= 16'd23487);
assign fi_addres[1353] = valid_point & (angle > 16'd23487 & angle <= 16'd23505);
assign fi_addres[1354] = valid_point & (angle > 16'd23505 & angle <= 16'd23523);
assign fi_addres[1355] = valid_point & (angle > 16'd23523 & angle <= 16'd23532);
assign fi_addres[1356] = valid_point & (angle > 16'd23532 & angle <= 16'd23550);
assign fi_addres[1357] = valid_point & (angle > 16'd23550 & angle <= 16'd23568);
assign fi_addres[1358] = valid_point & (angle > 16'd23568 & angle <= 16'd23586);
assign fi_addres[1359] = valid_point & (angle > 16'd23586 & angle <= 16'd23604);
assign fi_addres[1360] = valid_point & (angle > 16'd23604 & angle <= 16'd23622);
assign fi_addres[1361] = valid_point & (angle > 16'd23622 & angle <= 16'd23631);
assign fi_addres[1362] = valid_point & (angle > 16'd23631 & angle <= 16'd23649);
assign fi_addres[1363] = valid_point & (angle > 16'd23649 & angle <= 16'd23667);
assign fi_addres[1364] = valid_point & (angle > 16'd23667 & angle <= 16'd23685);
assign fi_addres[1365] = valid_point & (angle > 16'd23685 & angle <= 16'd23703);
assign fi_addres[1366] = valid_point & (angle > 16'd23703 & angle <= 16'd23721);
assign fi_addres[1367] = valid_point & (angle > 16'd23721 & angle <= 16'd23739);
assign fi_addres[1368] = valid_point & (angle > 16'd23739 & angle <= 16'd23757);
assign fi_addres[1369] = valid_point & (angle > 16'd23757 & angle <= 16'd23766);
assign fi_addres[1370] = valid_point & (angle > 16'd23766 & angle <= 16'd23784);
assign fi_addres[1371] = valid_point & (angle > 16'd23784 & angle <= 16'd23802);
assign fi_addres[1372] = valid_point & (angle > 16'd23802 & angle <= 16'd23820);
assign fi_addres[1373] = valid_point & (angle > 16'd23820 & angle <= 16'd23838);
assign fi_addres[1374] = valid_point & (angle > 16'd23838 & angle <= 16'd23855);
assign fi_addres[1375] = valid_point & (angle > 16'd23855 & angle <= 16'd23874);
assign fi_addres[1376] = valid_point & (angle > 16'd23874 & angle <= 16'd23882);
assign fi_addres[1377] = valid_point & (angle > 16'd23882 & angle <= 16'd23901);
assign fi_addres[1378] = valid_point & (angle > 16'd23901 & angle <= 16'd23919);
assign fi_addres[1379] = valid_point & (angle > 16'd23919 & angle <= 16'd23936);
assign fi_addres[1380] = valid_point & (angle > 16'd23936 & angle <= 16'd23955);
assign fi_addres[1381] = valid_point & (angle > 16'd23955 & angle <= 16'd23973);
assign fi_addres[1382] = valid_point & (angle > 16'd23973 & angle <= 16'd23991);
assign fi_addres[1383] = valid_point & (angle > 16'd23991 & angle <= 16'd23999);
assign fi_addres[1384] = valid_point & (angle > 16'd23999 & angle <= 16'd24017);
assign fi_addres[1385] = valid_point & (angle > 16'd24017 & angle <= 16'd24036);
assign fi_addres[1386] = valid_point & (angle > 16'd24036 & angle <= 16'd24054);
assign fi_addres[1387] = valid_point & (angle > 16'd24054 & angle <= 16'd24071);
assign fi_addres[1388] = valid_point & (angle > 16'd24071 & angle <= 16'd24089);
assign fi_addres[1389] = valid_point & (angle > 16'd24089 & angle <= 16'd24107);
assign fi_addres[1390] = valid_point & (angle > 16'd24107 & angle <= 16'd24116);
assign fi_addres[1391] = valid_point & (angle > 16'd24116 & angle <= 16'd24134);
assign fi_addres[1392] = valid_point & (angle > 16'd24134 & angle <= 16'd24152);
assign fi_addres[1393] = valid_point & (angle > 16'd24152 & angle <= 16'd24170);
assign fi_addres[1394] = valid_point & (angle > 16'd24170 & angle <= 16'd24188);
assign fi_addres[1395] = valid_point & (angle > 16'd24188 & angle <= 16'd24206);
assign fi_addres[1396] = valid_point & (angle > 16'd24206 & angle <= 16'd24224);
assign fi_addres[1397] = valid_point & (angle > 16'd24224 & angle <= 16'd24242);
assign fi_addres[1398] = valid_point & (angle > 16'd24242 & angle <= 16'd24251);
assign fi_addres[1399] = valid_point & (angle > 16'd24251 & angle <= 16'd24269);
assign fi_addres[1400] = valid_point & (angle > 16'd24269 & angle <= 16'd24287);
assign fi_addres[1401] = valid_point & (angle > 16'd24287 & angle <= 16'd24305);
assign fi_addres[1402] = valid_point & (angle > 16'd24305 & angle <= 16'd24323);
assign fi_addres[1403] = valid_point & (angle > 16'd24323 & angle <= 16'd24341);
assign fi_addres[1404] = valid_point & (angle > 16'd24341 & angle <= 16'd24359);
assign fi_addres[1405] = valid_point & (angle > 16'd24359 & angle <= 16'd24368);
assign fi_addres[1406] = valid_point & (angle > 16'd24368 & angle <= 16'd24386);
assign fi_addres[1407] = valid_point & (angle > 16'd24386 & angle <= 16'd24404);
assign fi_addres[1408] = valid_point & (angle > 16'd24404 & angle <= 16'd24422);
assign fi_addres[1409] = valid_point & (angle > 16'd24422 & angle <= 16'd24440);
assign fi_addres[1410] = valid_point & (angle > 16'd24440 & angle <= 16'd24458);
assign fi_addres[1411] = valid_point & (angle > 16'd24458 & angle <= 16'd24476);
assign fi_addres[1412] = valid_point & (angle > 16'd24476 & angle <= 16'd24494);
assign fi_addres[1413] = valid_point & (angle > 16'd24494 & angle <= 16'd24503);
assign fi_addres[1414] = valid_point & (angle > 16'd24503 & angle <= 16'd24521);
assign fi_addres[1415] = valid_point & (angle > 16'd24521 & angle <= 16'd24539);
assign fi_addres[1416] = valid_point & (angle > 16'd24539 & angle <= 16'd24557);
assign fi_addres[1417] = valid_point & (angle > 16'd24557 & angle <= 16'd24575);
assign fi_addres[1418] = valid_point & (angle > 16'd24575 & angle <= 16'd24593);
assign fi_addres[1419] = valid_point & (angle > 16'd24593 & angle <= 16'd24611);
assign fi_addres[1420] = valid_point & (angle > 16'd24611 & angle <= 16'd24620);
assign fi_addres[1421] = valid_point & (angle > 16'd24620 & angle <= 16'd24638);
assign fi_addres[1422] = valid_point & (angle > 16'd24638 & angle <= 16'd24656);
assign fi_addres[1423] = valid_point & (angle > 16'd24656 & angle <= 16'd24674);
assign fi_addres[1424] = valid_point & (angle > 16'd24674 & angle <= 16'd24692);
assign fi_addres[1425] = valid_point & (angle > 16'd24692 & angle <= 16'd24710);
assign fi_addres[1426] = valid_point & (angle > 16'd24710 & angle <= 16'd24728);
assign fi_addres[1427] = valid_point & (angle > 16'd24728 & angle <= 16'd24737);
assign fi_addres[1428] = valid_point & (angle > 16'd24737 & angle <= 16'd24755);
assign fi_addres[1429] = valid_point & (angle > 16'd24755 & angle <= 16'd24773);
assign fi_addres[1430] = valid_point & (angle > 16'd24773 & angle <= 16'd24791);
assign fi_addres[1431] = valid_point & (angle > 16'd24791 & angle <= 16'd24809);
assign fi_addres[1432] = valid_point & (angle > 16'd24809 & angle <= 16'd24827);
assign fi_addres[1433] = valid_point & (angle > 16'd24827 & angle <= 16'd24845);
assign fi_addres[1434] = valid_point & (angle > 16'd24845 & angle <= 16'd24854);
assign fi_addres[1435] = valid_point & (angle > 16'd24854 & angle <= 16'd24872);
assign fi_addres[1436] = valid_point & (angle > 16'd24872 & angle <= 16'd24890);
assign fi_addres[1437] = valid_point & (angle > 16'd24890 & angle <= 16'd24908);
assign fi_addres[1438] = valid_point & (angle > 16'd24908 & angle <= 16'd24926);
assign fi_addres[1439] = valid_point & (angle > 16'd24926 & angle <= 16'd24944);
assign fi_addres[1440] = valid_point & (angle > 16'd24944 & angle <= 16'd24962);
assign fi_addres[1441] = valid_point & (angle > 16'd24962 & angle <= 16'd24971);
assign fi_addres[1442] = valid_point & (angle > 16'd24971 & angle <= 16'd24989);
assign fi_addres[1443] = valid_point & (angle > 16'd24989 & angle <= 16'd25007);
assign fi_addres[1444] = valid_point & (angle > 16'd25007 & angle <= 16'd25025);
assign fi_addres[1445] = valid_point & (angle > 16'd25025 & angle <= 16'd25043);
assign fi_addres[1446] = valid_point & (angle > 16'd25043 & angle <= 16'd25061);
assign fi_addres[1447] = valid_point & (angle > 16'd25061 & angle <= 16'd25079);
assign fi_addres[1448] = valid_point & (angle > 16'd25079 & angle <= 16'd25088);
assign fi_addres[1449] = valid_point & (angle > 16'd25088 & angle <= 16'd25106);
assign fi_addres[1450] = valid_point & (angle > 16'd25106 & angle <= 16'd25124);
assign fi_addres[1451] = valid_point & (angle > 16'd25124 & angle <= 16'd25142);
assign fi_addres[1452] = valid_point & (angle > 16'd25142 & angle <= 16'd25160);
assign fi_addres[1453] = valid_point & (angle > 16'd25160 & angle <= 16'd25178);
assign fi_addres[1454] = valid_point & (angle > 16'd25178 & angle <= 16'd25196);
assign fi_addres[1455] = valid_point & (angle > 16'd25196 & angle <= 16'd25214);
assign fi_addres[1456] = valid_point & (angle > 16'd25214 & angle <= 16'd25223);
assign fi_addres[1457] = valid_point & (angle > 16'd25223 & angle <= 16'd25241);
assign fi_addres[1458] = valid_point & (angle > 16'd25241 & angle <= 16'd25259);
assign fi_addres[1459] = valid_point & (angle > 16'd25259 & angle <= 16'd25277);
assign fi_addres[1460] = valid_point & (angle > 16'd25277 & angle <= 16'd25294);
assign fi_addres[1461] = valid_point & (angle > 16'd25294 & angle <= 16'd25313);
assign fi_addres[1462] = valid_point & (angle > 16'd25313 & angle <= 16'd25331);
assign fi_addres[1463] = valid_point & (angle > 16'd25331 & angle <= 16'd25339);
assign fi_addres[1464] = valid_point & (angle > 16'd25339 & angle <= 16'd25357);
assign fi_addres[1465] = valid_point & (angle > 16'd25357 & angle <= 16'd25376);
assign fi_addres[1466] = valid_point & (angle > 16'd25376 & angle <= 16'd25394);
assign fi_addres[1467] = valid_point & (angle > 16'd25394 & angle <= 16'd25411);
assign fi_addres[1468] = valid_point & (angle > 16'd25411 & angle <= 16'd25429);
assign fi_addres[1469] = valid_point & (angle > 16'd25429 & angle <= 16'd25447);
assign fi_addres[1470] = valid_point & (angle > 16'd25447 & angle <= 16'd25457);
assign fi_addres[1471] = valid_point & (angle > 16'd25457 & angle <= 16'd25474);
assign fi_addres[1472] = valid_point & (angle > 16'd25474 & angle <= 16'd25492);
assign fi_addres[1473] = valid_point & (angle > 16'd25492 & angle <= 16'd25511);
assign fi_addres[1474] = valid_point & (angle > 16'd25511 & angle <= 16'd25528);
assign fi_addres[1475] = valid_point & (angle > 16'd25528 & angle <= 16'd25546);
assign fi_addres[1476] = valid_point & (angle > 16'd25546 & angle <= 16'd25565);
assign fi_addres[1477] = valid_point & (angle > 16'd25565 & angle <= 16'd25574);
assign fi_addres[1478] = valid_point & (angle > 16'd25574 & angle <= 16'd25591);
assign fi_addres[1479] = valid_point & (angle > 16'd25591 & angle <= 16'd25609);
assign fi_addres[1480] = valid_point & (angle > 16'd25609 & angle <= 16'd25627);
assign fi_addres[1481] = valid_point & (angle > 16'd25627 & angle <= 16'd25645);
assign fi_addres[1482] = valid_point & (angle > 16'd25645 & angle <= 16'd25663);
assign fi_addres[1483] = valid_point & (angle > 16'd25663 & angle <= 16'd25682);
assign fi_addres[1484] = valid_point & (angle > 16'd25682 & angle <= 16'd25691);
assign fi_addres[1485] = valid_point & (angle > 16'd25691 & angle <= 16'd25708);
assign fi_addres[1486] = valid_point & (angle > 16'd25708 & angle <= 16'd25726);
assign fi_addres[1487] = valid_point & (angle > 16'd25726 & angle <= 16'd25744);
assign fi_addres[1488] = valid_point & (angle > 16'd25744 & angle <= 16'd25762);
assign fi_addres[1489] = valid_point & (angle > 16'd25762 & angle <= 16'd25780);
assign fi_addres[1490] = valid_point & (angle > 16'd25780 & angle <= 16'd25798);
assign fi_addres[1491] = valid_point & (angle > 16'd25798 & angle <= 16'd25816);
assign fi_addres[1492] = valid_point & (angle > 16'd25816 & angle <= 16'd25825);
assign fi_addres[1493] = valid_point & (angle > 16'd25825 & angle <= 16'd25843);
assign fi_addres[1494] = valid_point & (angle > 16'd25843 & angle <= 16'd25862);
assign fi_addres[1495] = valid_point & (angle > 16'd25862 & angle <= 16'd25879);
assign fi_addres[1496] = valid_point & (angle > 16'd25879 & angle <= 16'd25898);
assign fi_addres[1497] = valid_point & (angle > 16'd25898 & angle <= 16'd25915);
assign fi_addres[1498] = valid_point & (angle > 16'd25915 & angle <= 16'd25933);
assign fi_addres[1499] = valid_point & (angle > 16'd25933 & angle <= 16'd25942);
assign fi_addres[1500] = valid_point & (angle > 16'd25942 & angle <= 16'd25960);
assign fi_addres[1501] = valid_point & (angle > 16'd25960 & angle <= 16'd25978);
assign fi_addres[1502] = valid_point & (angle > 16'd25978 & angle <= 16'd25996);
assign fi_addres[1503] = valid_point & (angle > 16'd25996 & angle <= 16'd26014);
assign fi_addres[1504] = valid_point & (angle > 16'd26014 & angle <= 16'd26032);
assign fi_addres[1505] = valid_point & (angle > 16'd26032 & angle <= 16'd26050);
assign fi_addres[1506] = valid_point & (angle > 16'd26050 & angle <= 16'd26059);
assign fi_addres[1507] = valid_point & (angle > 16'd26059 & angle <= 16'd26078);
assign fi_addres[1508] = valid_point & (angle > 16'd26078 & angle <= 16'd26096);
assign fi_addres[1509] = valid_point & (angle > 16'd26096 & angle <= 16'd26114);
assign fi_addres[1510] = valid_point & (angle > 16'd26114 & angle <= 16'd26132);
assign fi_addres[1511] = valid_point & (angle > 16'd26132 & angle <= 16'd26149);
assign fi_addres[1512] = valid_point & (angle > 16'd26149 & angle <= 16'd26168);
assign fi_addres[1513] = valid_point & (angle > 16'd26168 & angle <= 16'd26185);
assign fi_addres[1514] = valid_point & (angle > 16'd26185 & angle <= 16'd26194);
assign fi_addres[1515] = valid_point & (angle > 16'd26194 & angle <= 16'd26212);
assign fi_addres[1516] = valid_point & (angle > 16'd26212 & angle <= 16'd26230);
assign fi_addres[1517] = valid_point & (angle > 16'd26230 & angle <= 16'd26249);
assign fi_addres[1518] = valid_point & (angle > 16'd26249 & angle <= 16'd26266);
assign fi_addres[1519] = valid_point & (angle > 16'd26266 & angle <= 16'd26285);
assign fi_addres[1520] = valid_point & (angle > 16'd26285 & angle <= 16'd26302);
assign fi_addres[1521] = valid_point & (angle > 16'd26302 & angle <= 16'd26311);
assign fi_addres[1522] = valid_point & (angle > 16'd26311 & angle <= 16'd26329);
assign fi_addres[1523] = valid_point & (angle > 16'd26329 & angle <= 16'd26348);
assign fi_addres[1524] = valid_point & (angle > 16'd26348 & angle <= 16'd26365);
assign fi_addres[1525] = valid_point & (angle > 16'd26365 & angle <= 16'd26383);
assign fi_addres[1526] = valid_point & (angle > 16'd26383 & angle <= 16'd26402);
assign fi_addres[1527] = valid_point & (angle > 16'd26402 & angle <= 16'd26420);
assign fi_addres[1528] = valid_point & (angle > 16'd26420 & angle <= 16'd26429);
assign fi_addres[1529] = valid_point & (angle > 16'd26429 & angle <= 16'd26446);
assign fi_addres[1530] = valid_point & (angle > 16'd26446 & angle <= 16'd26464);
assign fi_addres[1531] = valid_point & (angle > 16'd26464 & angle <= 16'd26482);
assign fi_addres[1532] = valid_point & (angle > 16'd26482 & angle <= 16'd26500);
assign fi_addres[1533] = valid_point & (angle > 16'd26500 & angle <= 16'd26518);
assign fi_addres[1534] = valid_point & (angle > 16'd26518 & angle <= 16'd26536);
assign fi_addres[1535] = valid_point & (angle > 16'd26536 & angle <= 16'd26545);
assign fi_addres[1536] = valid_point & (angle > 16'd26545 & angle <= 16'd26564);
assign fi_addres[1537] = valid_point & (angle > 16'd26564 & angle <= 16'd26581);
assign fi_addres[1538] = valid_point & (angle > 16'd26581 & angle <= 16'd26600);
assign fi_addres[1539] = valid_point & (angle > 16'd26600 & angle <= 16'd26618);
assign fi_addres[1540] = valid_point & (angle > 16'd26618 & angle <= 16'd26636);
assign fi_addres[1541] = valid_point & (angle > 16'd26636 & angle <= 16'd26653);
assign fi_addres[1542] = valid_point & (angle > 16'd26653 & angle <= 16'd26662);
assign fi_addres[1543] = valid_point & (angle > 16'd26662 & angle <= 16'd26681);
assign fi_addres[1544] = valid_point & (angle > 16'd26681 & angle <= 16'd26698);
assign fi_addres[1545] = valid_point & (angle > 16'd26698 & angle <= 16'd26716);
assign fi_addres[1546] = valid_point & (angle > 16'd26716 & angle <= 16'd26735);
assign fi_addres[1547] = valid_point & (angle > 16'd26735 & angle <= 16'd26752);
assign fi_addres[1548] = valid_point & (angle > 16'd26752 & angle <= 16'd26771);
assign fi_addres[1549] = valid_point & (angle > 16'd26771 & angle <= 16'd26788);
assign fi_addres[1550] = valid_point & (angle > 16'd26788 & angle <= 16'd26797);
assign fi_addres[1551] = valid_point & (angle > 16'd26797 & angle <= 16'd26815);
assign fi_addres[1552] = valid_point & (angle > 16'd26815 & angle <= 16'd26833);
assign fi_addres[1553] = valid_point & (angle > 16'd26833 & angle <= 16'd26851);
assign fi_addres[1554] = valid_point & (angle > 16'd26851 & angle <= 16'd26869);
assign fi_addres[1555] = valid_point & (angle > 16'd26869 & angle <= 16'd26887);
assign fi_addres[1556] = valid_point & (angle > 16'd26887 & angle <= 16'd26906);
assign fi_addres[1557] = valid_point & (angle > 16'd26906 & angle <= 16'd26914);
assign fi_addres[1558] = valid_point & (angle > 16'd26914 & angle <= 16'd26932);
assign fi_addres[1559] = valid_point & (angle > 16'd26932 & angle <= 16'd26950);
assign fi_addres[1560] = valid_point & (angle > 16'd26950 & angle <= 16'd26969);
assign fi_addres[1561] = valid_point & (angle > 16'd26969 & angle <= 16'd26987);
assign fi_addres[1562] = valid_point & (angle > 16'd26987 & angle <= 16'd27004);
assign fi_addres[1563] = valid_point & (angle > 16'd27004 & angle <= 16'd27022);
assign fi_addres[1564] = valid_point & (angle > 16'd27022 & angle <= 16'd27031);
assign fi_addres[1565] = valid_point & (angle > 16'd27031 & angle <= 16'd27049);
assign fi_addres[1566] = valid_point & (angle > 16'd27049 & angle <= 16'd27067);
assign fi_addres[1567] = valid_point & (angle > 16'd27067 & angle <= 16'd27085);
assign fi_addres[1568] = valid_point & (angle > 16'd27085 & angle <= 16'd27103);
assign fi_addres[1569] = valid_point & (angle > 16'd27103 & angle <= 16'd27121);
assign fi_addres[1570] = valid_point & (angle > 16'd27121 & angle <= 16'd27139);
assign fi_addres[1571] = valid_point & (angle > 16'd27139 & angle <= 16'd27148);
assign fi_addres[1572] = valid_point & (angle > 16'd27148 & angle <= 16'd27167);
assign fi_addres[1573] = valid_point & (angle > 16'd27167 & angle <= 16'd27184);
assign fi_addres[1574] = valid_point & (angle > 16'd27184 & angle <= 16'd27202);
assign fi_addres[1575] = valid_point & (angle > 16'd27202 & angle <= 16'd27220);
assign fi_addres[1576] = valid_point & (angle > 16'd27220 & angle <= 16'd27238);
assign fi_addres[1577] = valid_point & (angle > 16'd27238 & angle <= 16'd27256);
assign fi_addres[1578] = valid_point & (angle > 16'd27256 & angle <= 16'd27265);
assign fi_addres[1579] = valid_point & (angle > 16'd27265 & angle <= 16'd27283);
assign fi_addres[1580] = valid_point & (angle > 16'd27283 & angle <= 16'd27302);
assign fi_addres[1581] = valid_point & (angle > 16'd27302 & angle <= 16'd27319);
assign fi_addres[1582] = valid_point & (angle > 16'd27319 & angle <= 16'd27337);
assign fi_addres[1583] = valid_point & (angle > 16'd27337 & angle <= 16'd27355);
assign fi_addres[1584] = valid_point & (angle > 16'd27355 & angle <= 16'd27374);
assign fi_addres[1585] = valid_point & (angle > 16'd27374 & angle <= 16'd27382);
assign fi_addres[1586] = valid_point & (angle > 16'd27382 & angle <= 16'd27400);
assign fi_addres[1587] = valid_point & (angle > 16'd27400 & angle <= 16'd27418);
assign fi_addres[1588] = valid_point & (angle > 16'd27418 & angle <= 16'd27437);
assign fi_addres[1589] = valid_point & (angle > 16'd27437 & angle <= 16'd27454);
assign fi_addres[1590] = valid_point & (angle > 16'd27454 & angle <= 16'd27473);
assign fi_addres[1591] = valid_point & (angle > 16'd27473 & angle <= 16'd27491);
assign fi_addres[1592] = valid_point & (angle > 16'd27491 & angle <= 16'd27509);
assign fi_addres[1593] = valid_point & (angle > 16'd27509 & angle <= 16'd27518);
assign fi_addres[1594] = valid_point & (angle > 16'd27518 & angle <= 16'd27535);
assign fi_addres[1595] = valid_point & (angle > 16'd27535 & angle <= 16'd27553);
assign fi_addres[1596] = valid_point & (angle > 16'd27553 & angle <= 16'd27572);
assign fi_addres[1597] = valid_point & (angle > 16'd27572 & angle <= 16'd27589);
assign fi_addres[1598] = valid_point & (angle > 16'd27589 & angle <= 16'd27607);
assign fi_addres[1599] = valid_point & (angle > 16'd27607 & angle <= 16'd27626);
assign fi_addres[1600] = valid_point & (angle > 16'd27626 & angle <= 16'd27634);
assign fi_addres[1601] = valid_point & (angle > 16'd27634 & angle <= 16'd27652);
assign fi_addres[1602] = valid_point & (angle > 16'd27652 & angle <= 16'd27671);
assign fi_addres[1603] = valid_point & (angle > 16'd27671 & angle <= 16'd27688);
assign fi_addres[1604] = valid_point & (angle > 16'd27688 & angle <= 16'd27707);
assign fi_addres[1605] = valid_point & (angle > 16'd27707 & angle <= 16'd27725);
assign fi_addres[1606] = valid_point & (angle > 16'd27725 & angle <= 16'd27742);
assign fi_addres[1607] = valid_point & (angle > 16'd27742 & angle <= 16'd27751);
assign fi_addres[1608] = valid_point & (angle > 16'd27751 & angle <= 16'd27770);
assign fi_addres[1609] = valid_point & (angle > 16'd27770 & angle <= 16'd27788);
assign fi_addres[1610] = valid_point & (angle > 16'd27788 & angle <= 16'd27806);
assign fi_addres[1611] = valid_point & (angle > 16'd27806 & angle <= 16'd27824);
assign fi_addres[1612] = valid_point & (angle > 16'd27824 & angle <= 16'd27842);
assign fi_addres[1613] = valid_point & (angle > 16'd27842 & angle <= 16'd27860);
assign fi_addres[1614] = valid_point & (angle > 16'd27860 & angle <= 16'd27869);
assign fi_addres[1615] = valid_point & (angle > 16'd27869 & angle <= 16'd27887);
assign fi_addres[1616] = valid_point & (angle > 16'd27887 & angle <= 16'd27905);
assign fi_addres[1617] = valid_point & (angle > 16'd27905 & angle <= 16'd27923);
assign fi_addres[1618] = valid_point & (angle > 16'd27923 & angle <= 16'd27941);
assign fi_addres[1619] = valid_point & (angle > 16'd27941 & angle <= 16'd27959);
assign fi_addres[1620] = valid_point & (angle > 16'd27959 & angle <= 16'd27977);
assign fi_addres[1621] = valid_point & (angle > 16'd27977 & angle <= 16'd27986);
assign fi_addres[1622] = valid_point & (angle > 16'd27986 & angle <= 16'd28004);
assign fi_addres[1623] = valid_point & (angle > 16'd28004 & angle <= 16'd28022);
assign fi_addres[1624] = valid_point & (angle > 16'd28022 & angle <= 16'd28040);
assign fi_addres[1625] = valid_point & (angle > 16'd28040 & angle <= 16'd28058);
assign fi_addres[1626] = valid_point & (angle > 16'd28058 & angle <= 16'd28076);
assign fi_addres[1627] = valid_point & (angle > 16'd28076 & angle <= 16'd28094);
assign fi_addres[1628] = valid_point & (angle > 16'd28094 & angle <= 16'd28112);
assign fi_addres[1629] = valid_point & (angle > 16'd28112 & angle <= 16'd28121);
assign fi_addres[1630] = valid_point & (angle > 16'd28121 & angle <= 16'd28139);
assign fi_addres[1631] = valid_point & (angle > 16'd28139 & angle <= 16'd28157);
assign fi_addres[1632] = valid_point & (angle > 16'd28157 & angle <= 16'd28175);
assign fi_addres[1633] = valid_point & (angle > 16'd28175 & angle <= 16'd28193);
assign fi_addres[1634] = valid_point & (angle > 16'd28193 & angle <= 16'd28210);
assign fi_addres[1635] = valid_point & (angle > 16'd28210 & angle <= 16'd28229);
assign fi_addres[1636] = valid_point & (angle > 16'd28229 & angle <= 16'd28237);
assign fi_addres[1637] = valid_point & (angle > 16'd28237 & angle <= 16'd28256);
assign fi_addres[1638] = valid_point & (angle > 16'd28256 & angle <= 16'd28274);
assign fi_addres[1639] = valid_point & (angle > 16'd28274 & angle <= 16'd28292);
assign fi_addres[1640] = valid_point & (angle > 16'd28292 & angle <= 16'd28310);
assign fi_addres[1641] = valid_point & (angle > 16'd28310 & angle <= 16'd28328);
assign fi_addres[1642] = valid_point & (angle > 16'd28328 & angle <= 16'd28346);
assign fi_addres[1643] = valid_point & (angle > 16'd28346 & angle <= 16'd28355);
assign fi_addres[1644] = valid_point & (angle > 16'd28355 & angle <= 16'd28373);
assign fi_addres[1645] = valid_point & (angle > 16'd28373 & angle <= 16'd28391);
assign fi_addres[1646] = valid_point & (angle > 16'd28391 & angle <= 16'd28409);
assign fi_addres[1647] = valid_point & (angle > 16'd28409 & angle <= 16'd28427);
assign fi_addres[1648] = valid_point & (angle > 16'd28427 & angle <= 16'd28445);
assign fi_addres[1649] = valid_point & (angle > 16'd28445 & angle <= 16'd28463);
assign fi_addres[1650] = valid_point & (angle > 16'd28463 & angle <= 16'd28472);
assign fi_addres[1651] = valid_point & (angle > 16'd28472 & angle <= 16'd28490);
assign fi_addres[1652] = valid_point & (angle > 16'd28490 & angle <= 16'd28508);
assign fi_addres[1653] = valid_point & (angle > 16'd28508 & angle <= 16'd28526);
assign fi_addres[1654] = valid_point & (angle > 16'd28526 & angle <= 16'd28544);
assign fi_addres[1655] = valid_point & (angle > 16'd28544 & angle <= 16'd28562);
assign fi_addres[1656] = valid_point & (angle > 16'd28562 & angle <= 16'd28580);
assign fi_addres[1657] = valid_point & (angle > 16'd28580 & angle <= 16'd28598);
assign fi_addres[1658] = valid_point & (angle > 16'd28598 & angle <= 16'd28607);
assign fi_addres[1659] = valid_point & (angle > 16'd28607 & angle <= 16'd28625);
assign fi_addres[1660] = valid_point & (angle > 16'd28625 & angle <= 16'd28643);
assign fi_addres[1661] = valid_point & (angle > 16'd28643 & angle <= 16'd28661);
assign fi_addres[1662] = valid_point & (angle > 16'd28661 & angle <= 16'd28679);
assign fi_addres[1663] = valid_point & (angle > 16'd28679 & angle <= 16'd28697);
assign fi_addres[1664] = valid_point & (angle > 16'd28697 & angle <= 16'd28715);
assign fi_addres[1665] = valid_point & (angle > 16'd28715 & angle <= 16'd28719);
assign fi_addres[1666] = valid_point & (angle > 16'd28719 & angle <= 16'd28742);
assign fi_addres[1667] = valid_point & (angle > 16'd28742 & angle <= 16'd28760);
assign fi_addres[1668] = valid_point & (angle > 16'd28760 & angle <= 16'd28772);
assign fi_addres[1669] = valid_point & (angle > 16'd28772 & angle <= 16'd28791);
assign fi_addres[1670] = valid_point & (angle > 16'd28791 & angle <= 16'd28809);
assign fi_addres[1671] = valid_point & (angle > 16'd28809 & angle <= 16'd28827);
assign fi_addres[1672] = valid_point & (angle > 16'd28827 & angle <= 16'd28836);
assign fi_addres[1673] = valid_point & (angle > 16'd28836 & angle <= 16'd28854);
assign fi_addres[1674] = valid_point & (angle > 16'd28854 & angle <= 16'd28872);
assign fi_addres[1675] = valid_point & (angle > 16'd28872 & angle <= 16'd28890);
assign fi_addres[1676] = valid_point & (angle > 16'd28890 & angle <= 16'd28907);
assign fi_addres[1677] = valid_point & (angle > 16'd28907 & angle <= 16'd28926);
assign fi_addres[1678] = valid_point & (angle > 16'd28926 & angle <= 16'd28943);
assign fi_addres[1679] = valid_point & (angle > 16'd28943 & angle <= 16'd28953);
assign fi_addres[1680] = valid_point & (angle > 16'd28953 & angle <= 16'd28971);
assign fi_addres[1681] = valid_point & (angle > 16'd28971 & angle <= 16'd28989);
assign fi_addres[1682] = valid_point & (angle > 16'd28989 & angle <= 16'd29007);
assign fi_addres[1683] = valid_point & (angle > 16'd29007 & angle <= 16'd29025);
assign fi_addres[1684] = valid_point & (angle > 16'd29025 & angle <= 16'd29048);
assign fi_addres[1685] = valid_point & (angle > 16'd29048 & angle <= 16'd29060);
assign fi_addres[1686] = valid_point & (angle > 16'd29060 & angle <= 16'd29070);
assign fi_addres[1687] = valid_point & (angle > 16'd29070 & angle <= 16'd29087);
assign fi_addres[1688] = valid_point & (angle > 16'd29087 & angle <= 16'd29105);
assign fi_addres[1689] = valid_point & (angle > 16'd29105 & angle <= 16'd29124);
assign fi_addres[1690] = valid_point & (angle > 16'd29124 & angle <= 16'd29141);
assign fi_addres[1691] = valid_point & (angle > 16'd29141 & angle <= 16'd29160);
assign fi_addres[1692] = valid_point & (angle > 16'd29160 & angle <= 16'd29177);
assign fi_addres[1693] = valid_point & (angle > 16'd29177 & angle <= 16'd29192);
assign fi_addres[1694] = valid_point & (angle > 16'd29192 & angle <= 16'd29210);
assign fi_addres[1695] = valid_point & (angle > 16'd29210 & angle <= 16'd29229);
assign fi_addres[1696] = valid_point & (angle > 16'd29229 & angle <= 16'd29246);
assign fi_addres[1697] = valid_point & (angle > 16'd29246 & angle <= 16'd29265);
assign fi_addres[1698] = valid_point & (angle > 16'd29265 & angle <= 16'd29283);
assign fi_addres[1699] = valid_point & (angle > 16'd29283 & angle <= 16'd29300);
assign fi_addres[1700] = valid_point & (angle > 16'd29300 & angle <= 16'd29310);
assign fi_addres[1701] = valid_point & (angle > 16'd29310 & angle <= 16'd29328);
assign fi_addres[1702] = valid_point & (angle > 16'd29328 & angle <= 16'd29346);
assign fi_addres[1703] = valid_point & (angle > 16'd29346 & angle <= 16'd29364);
assign fi_addres[1704] = valid_point & (angle > 16'd29364 & angle <= 16'd29382);
assign fi_addres[1705] = valid_point & (angle > 16'd29382 & angle <= 16'd29399);
assign fi_addres[1706] = valid_point & (angle > 16'd29399 & angle <= 16'd29418);
assign fi_addres[1707] = valid_point & (angle > 16'd29418 & angle <= 16'd29436);
assign fi_addres[1708] = valid_point & (angle > 16'd29436 & angle <= 16'd29445);
assign fi_addres[1709] = valid_point & (angle > 16'd29445 & angle <= 16'd29463);
assign fi_addres[1710] = valid_point & (angle > 16'd29463 & angle <= 16'd29475);
assign fi_addres[1711] = valid_point & (angle > 16'd29475 & angle <= 16'd29499);
assign fi_addres[1712] = valid_point & (angle > 16'd29499 & angle <= 16'd29511);
assign fi_addres[1713] = valid_point & (angle > 16'd29511 & angle <= 16'd29528);
assign fi_addres[1714] = valid_point & (angle > 16'd29528 & angle <= 16'd29553);
assign fi_addres[1715] = valid_point & (angle > 16'd29553 & angle <= 16'd29562);
assign fi_addres[1716] = valid_point & (angle > 16'd29562 & angle <= 16'd29580);
assign fi_addres[1717] = valid_point & (angle > 16'd29580 & angle <= 16'd29598);
assign fi_addres[1718] = valid_point & (angle > 16'd29598 & angle <= 16'd29616);
assign fi_addres[1719] = valid_point & (angle > 16'd29616 & angle <= 16'd29634);
assign fi_addres[1720] = valid_point & (angle > 16'd29634 & angle <= 16'd29652);
assign fi_addres[1721] = valid_point & (angle > 16'd29652 & angle <= 16'd29670);
assign fi_addres[1722] = valid_point & (angle > 16'd29670 & angle <= 16'd29679);
assign fi_addres[1723] = valid_point & (angle > 16'd29679 & angle <= 16'd29697);
assign fi_addres[1724] = valid_point & (angle > 16'd29697 & angle <= 16'd29715);
assign fi_addres[1725] = valid_point & (angle > 16'd29715 & angle <= 16'd29733);
assign fi_addres[1726] = valid_point & (angle > 16'd29733 & angle <= 16'd29751);
assign fi_addres[1727] = valid_point & (angle > 16'd29751 & angle <= 16'd29769);
assign fi_addres[1728] = valid_point & (angle > 16'd29769 & angle <= 16'd29782);
assign fi_addres[1729] = valid_point & (angle > 16'd29782 & angle <= 16'd29796);
assign fi_addres[1730] = valid_point & (angle > 16'd29796 & angle <= 16'd29810);
assign fi_addres[1731] = valid_point & (angle > 16'd29810 & angle <= 16'd29827);
assign fi_addres[1732] = valid_point & (angle > 16'd29827 & angle <= 16'd29845);
assign fi_addres[1733] = valid_point & (angle > 16'd29845 & angle <= 16'd29863);
assign fi_addres[1734] = valid_point & (angle > 16'd29863 & angle <= 16'd29881);
assign fi_addres[1735] = valid_point & (angle > 16'd29881 & angle <= 16'd29898);
assign fi_addres[1736] = valid_point & (angle > 16'd29898 & angle <= 16'd29908);
assign fi_addres[1737] = valid_point & (angle > 16'd29908 & angle <= 16'd29926);
assign fi_addres[1738] = valid_point & (angle > 16'd29926 & angle <= 16'd29944);
assign fi_addres[1739] = valid_point & (angle > 16'd29944 & angle <= 16'd29962);
assign fi_addres[1740] = valid_point & (angle > 16'd29962 & angle <= 16'd29980);
assign fi_addres[1741] = valid_point & (angle > 16'd29980 & angle <= 16'd29998);
assign fi_addres[1742] = valid_point & (angle > 16'd29998 & angle <= 16'd30016);
assign fi_addres[1743] = valid_point & (angle > 16'd30016 & angle <= 16'd30034);
assign fi_addres[1744] = valid_point & (angle > 16'd30034 & angle <= 16'd30043);
assign fi_addres[1745] = valid_point & (angle > 16'd30043 & angle <= 16'd30061);
assign fi_addres[1746] = valid_point & (angle > 16'd30061 & angle <= 16'd30079);
assign fi_addres[1747] = valid_point & (angle > 16'd30079 & angle <= 16'd30097);
assign fi_addres[1748] = valid_point & (angle > 16'd30097 & angle <= 16'd30115);
assign fi_addres[1749] = valid_point & (angle > 16'd30115 & angle <= 16'd30133);
assign fi_addres[1750] = valid_point & (angle > 16'd30133 & angle <= 16'd30151);
assign fi_addres[1751] = valid_point & (angle > 16'd30151 & angle <= 16'd30160);
assign fi_addres[1752] = valid_point & (angle > 16'd30160 & angle <= 16'd30178);
assign fi_addres[1753] = valid_point & (angle > 16'd30178 & angle <= 16'd30196);
assign fi_addres[1754] = valid_point & (angle > 16'd30196 & angle <= 16'd30214);
assign fi_addres[1755] = valid_point & (angle > 16'd30214 & angle <= 16'd30232);
assign fi_addres[1756] = valid_point & (angle > 16'd30232 & angle <= 16'd30250);
assign fi_addres[1757] = valid_point & (angle > 16'd30250 & angle <= 16'd30268);
assign fi_addres[1758] = valid_point & (angle > 16'd30268 & angle <= 16'd30277);
assign fi_addres[1759] = valid_point & (angle > 16'd30277 & angle <= 16'd30295);
assign fi_addres[1760] = valid_point & (angle > 16'd30295 & angle <= 16'd30313);
assign fi_addres[1761] = valid_point & (angle > 16'd30313 & angle <= 16'd30331);
assign fi_addres[1762] = valid_point & (angle > 16'd30331 & angle <= 16'd30349);
assign fi_addres[1763] = valid_point & (angle > 16'd30349 & angle <= 16'd30372);
assign fi_addres[1764] = valid_point & (angle > 16'd30372 & angle <= 16'd30385);
assign fi_addres[1765] = valid_point & (angle > 16'd30385 & angle <= 16'd30394);
assign fi_addres[1766] = valid_point & (angle > 16'd30394 & angle <= 16'd30412);
assign fi_addres[1767] = valid_point & (angle > 16'd30412 & angle <= 16'd30430);
assign fi_addres[1768] = valid_point & (angle > 16'd30430 & angle <= 16'd30448);
assign fi_addres[1769] = valid_point & (angle > 16'd30448 & angle <= 16'd30466);
assign fi_addres[1770] = valid_point & (angle > 16'd30466 & angle <= 16'd30484);
assign fi_addres[1771] = valid_point & (angle > 16'd30484 & angle <= 16'd30502);
assign fi_addres[1772] = valid_point & (angle > 16'd30502 & angle <= 16'd30511);
assign fi_addres[1773] = valid_point & (angle > 16'd30511 & angle <= 16'd30529);
assign fi_addres[1774] = valid_point & (angle > 16'd30529 & angle <= 16'd30547);
assign fi_addres[1775] = valid_point & (angle > 16'd30547 & angle <= 16'd30565);
assign fi_addres[1776] = valid_point & (angle > 16'd30565 & angle <= 16'd30582);
assign fi_addres[1777] = valid_point & (angle > 16'd30582 & angle <= 16'd30601);
assign fi_addres[1778] = valid_point & (angle > 16'd30601 & angle <= 16'd30625);
assign fi_addres[1779] = valid_point & (angle > 16'd30625 & angle <= 16'd30643);
assign fi_addres[1780] = valid_point & (angle > 16'd30643 & angle <= 16'd30652);
assign fi_addres[1781] = valid_point & (angle > 16'd30652 & angle <= 16'd30670);
assign fi_addres[1782] = valid_point & (angle > 16'd30670 & angle <= 16'd30688);
assign fi_addres[1783] = valid_point & (angle > 16'd30688 & angle <= 16'd30706);
assign fi_addres[1784] = valid_point & (angle > 16'd30706 & angle <= 16'd30724);
assign fi_addres[1785] = valid_point & (angle > 16'd30724 & angle <= 16'd30742);
assign fi_addres[1786] = valid_point & (angle > 16'd30742 & angle <= 16'd30760);
assign fi_addres[1787] = valid_point & (angle > 16'd30760 & angle <= 16'd30769);
assign fi_addres[1788] = valid_point & (angle > 16'd30769 & angle <= 16'd30787);
assign fi_addres[1789] = valid_point & (angle > 16'd30787 & angle <= 16'd30805);
assign fi_addres[1790] = valid_point & (angle > 16'd30805 & angle <= 16'd30823);
assign fi_addres[1791] = valid_point & (angle > 16'd30823 & angle <= 16'd30841);
assign fi_addres[1792] = valid_point & (angle > 16'd30841 & angle <= 16'd30859);
assign fi_addres[1793] = valid_point & (angle > 16'd30859 & angle <= 16'd30868);
assign fi_addres[1794] = valid_point & (angle > 16'd30868 & angle <= 16'd30886);
assign fi_addres[1795] = valid_point & (angle > 16'd30886 & angle <= 16'd30904);
assign fi_addres[1796] = valid_point & (angle > 16'd30904 & angle <= 16'd30922);
assign fi_addres[1797] = valid_point & (angle > 16'd30922 & angle <= 16'd30940);
assign fi_addres[1798] = valid_point & (angle > 16'd30940 & angle <= 16'd30958);
assign fi_addres[1799] = valid_point & (angle > 16'd30958 & angle <= 16'd30976);
assign fi_addres[1800] = valid_point & (angle > 16'd30976 & angle <= 16'd30994);
assign fi_addres[1801] = valid_point & (angle > 16'd30994 & angle <= 16'd31003);
assign fi_addres[1802] = valid_point & (angle > 16'd31003 & angle <= 16'd31021);
assign fi_addres[1803] = valid_point & (angle > 16'd31021 & angle <= 16'd31039);
assign fi_addres[1804] = valid_point & (angle > 16'd31039 & angle <= 16'd31057);
assign fi_addres[1805] = valid_point & (angle > 16'd31057 & angle <= 16'd31075);
assign fi_addres[1806] = valid_point & (angle > 16'd31075 & angle <= 16'd31093);
assign fi_addres[1807] = valid_point & (angle > 16'd31093 & angle <= 16'd31111);
assign fi_addres[1808] = valid_point & (angle > 16'd31111 & angle <= 16'd31120);
assign fi_addres[1809] = valid_point & (angle > 16'd31120 & angle <= 16'd31138);
assign fi_addres[1810] = valid_point & (angle > 16'd31138 & angle <= 16'd31156);
assign fi_addres[1811] = valid_point & (angle > 16'd31156 & angle <= 16'd31174);
assign fi_addres[1812] = valid_point & (angle > 16'd31174 & angle <= 16'd31192);
assign fi_addres[1813] = valid_point & (angle > 16'd31192 & angle <= 16'd31210);
assign fi_addres[1814] = valid_point & (angle > 16'd31210 & angle <= 16'd31228);
assign fi_addres[1815] = valid_point & (angle > 16'd31228 & angle <= 16'd31237);
assign fi_addres[1816] = valid_point & (angle > 16'd31237 & angle <= 16'd31255);
assign fi_addres[1817] = valid_point & (angle > 16'd31255 & angle <= 16'd31273);
assign fi_addres[1818] = valid_point & (angle > 16'd31273 & angle <= 16'd31291);
assign fi_addres[1819] = valid_point & (angle > 16'd31291 & angle <= 16'd31310);
assign fi_addres[1820] = valid_point & (angle > 16'd31310 & angle <= 16'd31328);
assign fi_addres[1821] = valid_point & (angle > 16'd31328 & angle <= 16'd31345);
assign fi_addres[1822] = valid_point & (angle > 16'd31345 & angle <= 16'd31354);
assign fi_addres[1823] = valid_point & (angle > 16'd31354 & angle <= 16'd31373);
assign fi_addres[1824] = valid_point & (angle > 16'd31373 & angle <= 16'd31391);
assign fi_addres[1825] = valid_point & (angle > 16'd31391 & angle <= 16'd31409);
assign fi_addres[1826] = valid_point & (angle > 16'd31409 & angle <= 16'd31423);
assign fi_addres[1827] = valid_point & (angle > 16'd31423 & angle <= 16'd31441);
assign fi_addres[1828] = valid_point & (angle > 16'd31441 & angle <= 16'd31459);
assign fi_addres[1829] = valid_point & (angle > 16'd31459 & angle <= 16'd31468);
assign fi_addres[1830] = valid_point & (angle > 16'd31468 & angle <= 16'd31486);
assign fi_addres[1831] = valid_point & (angle > 16'd31486 & angle <= 16'd31504);
assign fi_addres[1832] = valid_point & (angle > 16'd31504 & angle <= 16'd31522);
assign fi_addres[1833] = valid_point & (angle > 16'd31522 & angle <= 16'd31544);
assign fi_addres[1834] = valid_point & (angle > 16'd31544 & angle <= 16'd31558);
assign fi_addres[1835] = valid_point & (angle > 16'd31558 & angle <= 16'd31576);
assign fi_addres[1836] = valid_point & (angle > 16'd31576 & angle <= 16'd31594);
assign fi_addres[1837] = valid_point & (angle > 16'd31594 & angle <= 16'd31603);
assign fi_addres[1838] = valid_point & (angle > 16'd31603 & angle <= 16'd31621);
assign fi_addres[1839] = valid_point & (angle > 16'd31621 & angle <= 16'd31643);
assign fi_addres[1840] = valid_point & (angle > 16'd31643 & angle <= 16'd31661);
assign fi_addres[1841] = valid_point & (angle > 16'd31661 & angle <= 16'd31679);
assign fi_addres[1842] = valid_point & (angle > 16'd31679 & angle <= 16'd31697);
assign fi_addres[1843] = valid_point & (angle > 16'd31697 & angle <= 16'd31711);
assign fi_addres[1844] = valid_point & (angle > 16'd31711 & angle <= 16'd31720);
assign fi_addres[1845] = valid_point & (angle > 16'd31720 & angle <= 16'd31738);
assign fi_addres[1846] = valid_point & (angle > 16'd31738 & angle <= 16'd31756);
assign fi_addres[1847] = valid_point & (angle > 16'd31756 & angle <= 16'd31774);
assign fi_addres[1848] = valid_point & (angle > 16'd31774 & angle <= 16'd31792);
assign fi_addres[1849] = valid_point & (angle > 16'd31792 & angle <= 16'd31810);
assign fi_addres[1850] = valid_point & (angle > 16'd31810 & angle <= 16'd31828);
assign fi_addres[1851] = valid_point & (angle > 16'd31828 & angle <= 16'd31837);
assign fi_addres[1852] = valid_point & (angle > 16'd31837 & angle <= 16'd31855);
assign fi_addres[1853] = valid_point & (angle > 16'd31855 & angle <= 16'd31873);
assign fi_addres[1854] = valid_point & (angle > 16'd31873 & angle <= 16'd31891);
assign fi_addres[1855] = valid_point & (angle > 16'd31891 & angle <= 16'd31909);
assign fi_addres[1856] = valid_point & (angle > 16'd31909 & angle <= 16'd31927);
assign fi_addres[1857] = valid_point & (angle > 16'd31927 & angle <= 16'd31945);
assign fi_addres[1858] = valid_point & (angle > 16'd31945 & angle <= 16'd31958);
assign fi_addres[1859] = valid_point & (angle > 16'd31958 & angle <= 16'd31976);
assign fi_addres[1860] = valid_point & (angle > 16'd31976 & angle <= 16'd31994);
assign fi_addres[1861] = valid_point & (angle > 16'd31994 & angle <= 16'd32013);
assign fi_addres[1862] = valid_point & (angle > 16'd32013 & angle <= 16'd32026);
assign fi_addres[1863] = valid_point & (angle > 16'd32026 & angle <= 16'd32044);
assign fi_addres[1864] = valid_point & (angle > 16'd32044 & angle <= 16'd32062);
assign fi_addres[1865] = valid_point & (angle > 16'd32062 & angle <= 16'd32071);
assign fi_addres[1866] = valid_point & (angle > 16'd32071 & angle <= 16'd32089);
assign fi_addres[1867] = valid_point & (angle > 16'd32089 & angle <= 16'd32107);
assign fi_addres[1868] = valid_point & (angle > 16'd32107 & angle <= 16'd32125);
assign fi_addres[1869] = valid_point & (angle > 16'd32125 & angle <= 16'd32143);
assign fi_addres[1870] = valid_point & (angle > 16'd32143 & angle <= 16'd32161);
assign fi_addres[1871] = valid_point & (angle > 16'd32161 & angle <= 16'd32180);
assign fi_addres[1872] = valid_point & (angle > 16'd32180 & angle <= 16'd32189);
assign fi_addres[1873] = valid_point & (angle > 16'd32189 & angle <= 16'd32211);
assign fi_addres[1874] = valid_point & (angle > 16'd32211 & angle <= 16'd32229);
assign fi_addres[1875] = valid_point & (angle > 16'd32229 & angle <= 16'd32247);
assign fi_addres[1876] = valid_point & (angle > 16'd32247 & angle <= 16'd32265);
assign fi_addres[1877] = valid_point & (angle > 16'd32265 & angle <= 16'd32283);
assign fi_addres[1878] = valid_point & (angle > 16'd32283 & angle <= 16'd32301);
assign fi_addres[1879] = valid_point & (angle > 16'd32301 & angle <= 16'd32319);
assign fi_addres[1880] = valid_point & (angle > 16'd32319 & angle <= 16'd32328);
assign fi_addres[1881] = valid_point & (angle > 16'd32328 & angle <= 16'd32346);
assign fi_addres[1882] = valid_point & (angle > 16'd32346 & angle <= 16'd32364);
assign fi_addres[1883] = valid_point & (angle > 16'd32364 & angle <= 16'd32382);
assign fi_addres[1884] = valid_point & (angle > 16'd32382 & angle <= 16'd32400);
assign fi_addres[1885] = valid_point & (angle > 16'd32400 & angle <= 16'd32418);
assign fi_addres[1886] = valid_point & (angle > 16'd32418 & angle <= 16'd32436);
assign fi_addres[1887] = valid_point & (angle > 16'd32436 & angle <= 16'd32445);
assign fi_addres[1888] = valid_point & (angle > 16'd32445 & angle <= 16'd32463);
assign fi_addres[1889] = valid_point & (angle > 16'd32463 & angle <= 16'd32481);
assign fi_addres[1890] = valid_point & (angle > 16'd32481 & angle <= 16'd32499);
assign fi_addres[1891] = valid_point & (angle > 16'd32499 & angle <= 16'd32517);
assign fi_addres[1892] = valid_point & (angle > 16'd32517 & angle <= 16'd32535);
assign fi_addres[1893] = valid_point & (angle > 16'd32535 & angle <= 16'd32553);
assign fi_addres[1894] = valid_point & (angle > 16'd32553 & angle <= 16'd32562);
assign fi_addres[1895] = valid_point & (angle > 16'd32562 & angle <= 16'd32580);
assign fi_addres[1896] = valid_point & (angle > 16'd32580 & angle <= 16'd32598);
assign fi_addres[1897] = valid_point & (angle > 16'd32598 & angle <= 16'd32616);
assign fi_addres[1898] = valid_point & (angle > 16'd32616 & angle <= 16'd32634);
assign fi_addres[1899] = valid_point & (angle > 16'd32634 & angle <= 16'd32652);
assign fi_addres[1900] = valid_point & (angle > 16'd32652 & angle <= 16'd32670);
assign fi_addres[1901] = valid_point & (angle > 16'd32670 & angle <= 16'd32679);
assign fi_addres[1902] = valid_point & (angle > 16'd32679 & angle <= 16'd32697);
assign fi_addres[1903] = valid_point & (angle > 16'd32697 & angle <= 16'd32716);
assign fi_addres[1904] = valid_point & (angle > 16'd32716 & angle <= 16'd32733);
assign fi_addres[1905] = valid_point & (angle > 16'd32733 & angle <= 16'd32751);
assign fi_addres[1906] = valid_point & (angle > 16'd32751 & angle <= 16'd32769);
assign fi_addres[1907] = valid_point & (angle > 16'd32769 & angle <= 16'd32788);
assign fi_addres[1908] = valid_point & (angle > 16'd32788 & angle <= 16'd32797);
assign fi_addres[1909] = valid_point & (angle > 16'd32797 & angle <= 16'd32815);
assign fi_addres[1910] = valid_point & (angle > 16'd32815 & angle <= 16'd32833);
assign fi_addres[1911] = valid_point & (angle > 16'd32833 & angle <= 16'd32851);
assign fi_addres[1912] = valid_point & (angle > 16'd32851 & angle <= 16'd32869);
assign fi_addres[1913] = valid_point & (angle > 16'd32869 & angle <= 16'd32887);
assign fi_addres[1914] = valid_point & (angle > 16'd32887 & angle <= 16'd32905);
assign fi_addres[1915] = valid_point & (angle > 16'd32905 & angle <= 16'd32914);
assign fi_addres[1916] = valid_point & (angle > 16'd32914 & angle <= 16'd32932);
assign fi_addres[1917] = valid_point & (angle > 16'd32932 & angle <= 16'd32950);
assign fi_addres[1918] = valid_point & (angle > 16'd32950 & angle <= 16'd32968);
assign fi_addres[1919] = valid_point & (angle > 16'd32968 & angle <= 16'd32986);
assign fi_addres[1920] = valid_point & (angle > 16'd32986 & angle <= 16'd33004);
assign fi_addres[1921] = valid_point & (angle > 16'd33004 & angle <= 16'd33022);
assign fi_addres[1922] = valid_point & (angle > 16'd33022 & angle <= 16'd33040);
assign fi_addres[1923] = valid_point & (angle > 16'd33040 & angle <= 16'd33049);
assign fi_addres[1924] = valid_point & (angle > 16'd33049 & angle <= 16'd33067);
assign fi_addres[1925] = valid_point & (angle > 16'd33067 & angle <= 16'd33085);
assign fi_addres[1926] = valid_point & (angle > 16'd33085 & angle <= 16'd33103);
assign fi_addres[1927] = valid_point & (angle > 16'd33103 & angle <= 16'd33121);
assign fi_addres[1928] = valid_point & (angle > 16'd33121 & angle <= 16'd33139);
assign fi_addres[1929] = valid_point & (angle > 16'd33139 & angle <= 16'd33157);
assign fi_addres[1930] = valid_point & (angle > 16'd33157 & angle <= 16'd33166);
assign fi_addres[1931] = valid_point & (angle > 16'd33166 & angle <= 16'd33184);
assign fi_addres[1932] = valid_point & (angle > 16'd33184 & angle <= 16'd33202);
assign fi_addres[1933] = valid_point & (angle > 16'd33202 & angle <= 16'd33220);
assign fi_addres[1934] = valid_point & (angle > 16'd33220 & angle <= 16'd33238);
assign fi_addres[1935] = valid_point & (angle > 16'd33238 & angle <= 16'd33256);
assign fi_addres[1936] = valid_point & (angle > 16'd33256 & angle <= 16'd33274);
assign fi_addres[1937] = valid_point & (angle > 16'd33274 & angle <= 16'd33283);
assign fi_addres[1938] = valid_point & (angle > 16'd33283 & angle <= 16'd33301);
assign fi_addres[1939] = valid_point & (angle > 16'd33301 & angle <= 16'd33319);
assign fi_addres[1940] = valid_point & (angle > 16'd33319 & angle <= 16'd33337);
assign fi_addres[1941] = valid_point & (angle > 16'd33337 & angle <= 16'd33355);
assign fi_addres[1942] = valid_point & (angle > 16'd33355 & angle <= 16'd33374);
assign fi_addres[1943] = valid_point & (angle > 16'd33374 & angle <= 16'd33392);
assign fi_addres[1944] = valid_point & (angle > 16'd33392 & angle <= 16'd33401);
assign fi_addres[1945] = valid_point & (angle > 16'd33401 & angle <= 16'd33419);
assign fi_addres[1946] = valid_point & (angle > 16'd33419 & angle <= 16'd33437);
assign fi_addres[1947] = valid_point & (angle > 16'd33437 & angle <= 16'd33455);
assign fi_addres[1948] = valid_point & (angle > 16'd33455 & angle <= 16'd33473);
assign fi_addres[1949] = valid_point & (angle > 16'd33473 & angle <= 16'd33491);
assign fi_addres[1950] = valid_point & (angle > 16'd33491 & angle <= 16'd33509);
assign fi_addres[1951] = valid_point & (angle > 16'd33509 & angle <= 16'd33527);
assign fi_addres[1952] = valid_point & (angle > 16'd33527 & angle <= 16'd33554);
assign fi_addres[1953] = valid_point & (angle > 16'd33554 & angle <= 16'd33572);
assign fi_addres[1954] = valid_point & (angle > 16'd33572 & angle <= 16'd33590);
assign fi_addres[1955] = valid_point & (angle > 16'd33590 & angle <= 16'd33608);
assign fi_addres[1956] = valid_point & (angle > 16'd33608 & angle <= 16'd33626);
assign fi_addres[1957] = valid_point & (angle > 16'd33626 & angle <= 16'd33644);
assign fi_addres[1958] = valid_point & (angle > 16'd33644 & angle <= 16'd33654);
assign fi_addres[1959] = valid_point & (angle > 16'd33654 & angle <= 16'd33672);
assign fi_addres[1960] = valid_point & (angle > 16'd33672 & angle <= 16'd33689);
assign fi_addres[1961] = valid_point & (angle > 16'd33689 & angle <= 16'd33707);
assign fi_addres[1962] = valid_point & (angle > 16'd33707 & angle <= 16'd33725);
assign fi_addres[1963] = valid_point & (angle > 16'd33725 & angle <= 16'd33743);
assign fi_addres[1964] = valid_point & (angle > 16'd33743 & angle <= 16'd33761);
assign fi_addres[1965] = valid_point & (angle > 16'd33761 & angle <= 16'd33770);
assign fi_addres[1966] = valid_point & (angle > 16'd33770 & angle <= 16'd33788);
assign fi_addres[1967] = valid_point & (angle > 16'd33788 & angle <= 16'd33806);
assign fi_addres[1968] = valid_point & (angle > 16'd33806 & angle <= 16'd33824);
assign fi_addres[1969] = valid_point & (angle > 16'd33824 & angle <= 16'd33842);
assign fi_addres[1970] = valid_point & (angle > 16'd33842 & angle <= 16'd33860);
assign fi_addres[1971] = valid_point & (angle > 16'd33860 & angle <= 16'd33878);
assign fi_addres[1972] = valid_point & (angle > 16'd33878 & angle <= 16'd33887);
assign fi_addres[1973] = valid_point & (angle > 16'd33887 & angle <= 16'd33906);
assign fi_addres[1974] = valid_point & (angle > 16'd33906 & angle <= 16'd33922);
assign fi_addres[1975] = valid_point & (angle > 16'd33922 & angle <= 16'd33940);
assign fi_addres[1976] = valid_point & (angle > 16'd33940 & angle <= 16'd33958);
assign fi_addres[1977] = valid_point & (angle > 16'd33958 & angle <= 16'd33976);
assign fi_addres[1978] = valid_point & (angle > 16'd33976 & angle <= 16'd33994);
assign fi_addres[1979] = valid_point & (angle > 16'd33994 & angle <= 16'd34003);
assign fi_addres[1980] = valid_point & (angle > 16'd34003 & angle <= 16'd34021);
assign fi_addres[1981] = valid_point & (angle > 16'd34021 & angle <= 16'd34039);
assign fi_addres[1982] = valid_point & (angle > 16'd34039 & angle <= 16'd34057);
assign fi_addres[1983] = valid_point & (angle > 16'd34057 & angle <= 16'd34077);
assign fi_addres[1984] = valid_point & (angle > 16'd34077 & angle <= 16'd34093);
assign fi_addres[1985] = valid_point & (angle > 16'd34093 & angle <= 16'd34111);
assign fi_addres[1986] = valid_point & (angle > 16'd34111 & angle <= 16'd34120);
assign fi_addres[1987] = valid_point & (angle > 16'd34120 & angle <= 16'd34138);
assign fi_addres[1988] = valid_point & (angle > 16'd34138 & angle <= 16'd34156);
assign fi_addres[1989] = valid_point & (angle > 16'd34156 & angle <= 16'd34174);
assign fi_addres[1990] = valid_point & (angle > 16'd34174 & angle <= 16'd34193);
assign fi_addres[1991] = valid_point & (angle > 16'd34193 & angle <= 16'd34212);
assign fi_addres[1992] = valid_point & (angle > 16'd34212 & angle <= 16'd34230);
assign fi_addres[1993] = valid_point & (angle > 16'd34230 & angle <= 16'd34239);
assign fi_addres[1994] = valid_point & (angle > 16'd34239 & angle <= 16'd34256);
assign fi_addres[1995] = valid_point & (angle > 16'd34256 & angle <= 16'd34274);
assign fi_addres[1996] = valid_point & (angle > 16'd34274 & angle <= 16'd34292);
assign fi_addres[1997] = valid_point & (angle > 16'd34292 & angle <= 16'd34311);
assign fi_addres[1998] = valid_point & (angle > 16'd34311 & angle <= 16'd34329);
assign fi_addres[1999] = valid_point & (angle > 16'd34329 & angle <= 16'd34346);
assign fi_addres[2000] = valid_point & (angle > 16'd34346 & angle <= 16'd34364);
assign fi_addres[2001] = valid_point & (angle > 16'd34364 & angle <= 16'd34373);
assign fi_addres[2002] = valid_point & (angle > 16'd34373 & angle <= 16'd34391);
assign fi_addres[2003] = valid_point & (angle > 16'd34391 & angle <= 16'd34422);
assign fi_addres[2004] = valid_point & (angle > 16'd34422 & angle <= 16'd34445);
assign fi_addres[2005] = valid_point & (angle > 16'd34445 & angle <= 16'd34463);
assign fi_addres[2006] = valid_point & (angle > 16'd34463 & angle <= 16'd34481);
assign fi_addres[2007] = valid_point & (angle > 16'd34481 & angle <= 16'd34503);
assign fi_addres[2008] = valid_point & (angle > 16'd34503 & angle <= 16'd34521);
assign fi_addres[2009] = valid_point & (angle > 16'd34521 & angle <= 16'd34539);
assign fi_addres[2010] = valid_point & (angle > 16'd34539 & angle <= 16'd34566);
assign fi_addres[2011] = valid_point & (angle > 16'd34566 & angle <= 16'd34584);
assign fi_addres[2012] = valid_point & (angle > 16'd34584 & angle <= 16'd34607);
assign fi_addres[2013] = valid_point & (angle > 16'd34607 & angle <= 16'd34629);
assign fi_addres[2014] = valid_point & (angle > 16'd34629 & angle <= 16'd34647);
assign fi_addres[2015] = valid_point & (angle > 16'd34647 & angle <= 16'd34665);
assign fi_addres[2016] = valid_point & (angle > 16'd34665 & angle <= 16'd34696);
assign fi_addres[2017] = valid_point & (angle > 16'd34696 & angle <= 16'd34715);
assign fi_addres[2018] = valid_point & (angle > 16'd34715 & angle <= 16'd34732);
assign fi_addres[2019] = valid_point & (angle > 16'd34732 & angle <= 16'd34748);
assign fi_addres[2020] = valid_point & (angle > 16'd34748 & angle <= 16'd34773);
assign fi_addres[2021] = valid_point & (angle > 16'd34773 & angle <= 16'd34800);
assign fi_addres[2022] = valid_point & (angle > 16'd34800 & angle <= 16'd34818);
assign fi_addres[2023] = valid_point & (angle > 16'd34818 & angle <= 16'd34845);
assign fi_addres[2024] = valid_point & (angle > 16'd34845 & angle <= 16'd34863);
assign fi_addres[2025] = valid_point & (angle > 16'd34863 & angle <= 16'd34885);
assign fi_addres[2026] = valid_point & (angle > 16'd34885 & angle <= 16'd34903);
assign fi_addres[2027] = valid_point & (angle > 16'd34903 & angle <= 16'd34934);
assign fi_addres[2028] = valid_point & (angle > 16'd34934 & angle <= 16'd34952);
assign fi_addres[2029] = valid_point & (angle > 16'd34952 & angle <= 16'd34979);
assign fi_addres[2030] = valid_point & (angle > 16'd34979 & angle <= 16'd34995);
assign fi_addres[2031] = valid_point & (angle > 16'd34995 & angle <= 16'd35013);
assign fi_addres[2032] = valid_point & (angle > 16'd35013 & angle <= 16'd35031);
assign fi_addres[2033] = valid_point & (angle > 16'd35031 & angle <= 16'd35049);
assign fi_addres[2034] = valid_point & (angle > 16'd35049 & angle <= 16'd35067);
assign fi_addres[2035] = valid_point & (angle > 16'd35067 & angle <= 16'd35085);
assign fi_addres[2036] = valid_point & (angle > 16'd35085 & angle <= 16'd35094);
assign fi_addres[2037] = valid_point & (angle > 16'd35094 & angle <= 16'd35112);
assign fi_addres[2038] = valid_point & (angle > 16'd35112 & angle <= 16'd35133);
assign fi_addres[2039] = valid_point & (angle > 16'd35133 & angle <= 16'd35164);
assign fi_addres[2040] = valid_point & (angle > 16'd35164 & angle <= 16'd35182);
assign fi_addres[2041] = valid_point & (angle > 16'd35182 & angle <= 16'd35204);
assign fi_addres[2042] = valid_point & (angle > 16'd35204 & angle <= 16'd35227);
assign fi_addres[2043] = valid_point & (angle > 16'd35227 & angle <= 16'd35244);
assign fi_addres[2044] = valid_point & (angle > 16'd35244 & angle <= 16'd35263);
assign fi_addres[2045] = valid_point & (angle > 16'd35263 & angle <= 16'd35285);
assign fi_addres[2046] = valid_point & (angle > 16'd35285 & angle <= 16'd35303);
assign fi_addres[2047] = valid_point & (angle > 16'd35303 & angle <= 16'd35322);
assign fi_addres[2048] = valid_point & (angle > 16'd35322 & angle <= 16'd35343);
assign fi_addres[2049] = valid_point & (angle > 16'd35343 & angle <= 16'd35362);
assign fi_addres[2050] = valid_point & (angle > 16'd35362 & angle <= 16'd35385);
assign fi_addres[2051] = valid_point & (angle > 16'd35385 & angle <= 16'd35403);
assign fi_addres[2052] = valid_point & (angle > 16'd35403 & angle <= 16'd35421);
assign fi_addres[2053] = valid_point & (angle > 16'd35421 & angle <= 16'd35438);
assign fi_addres[2054] = valid_point & (angle > 16'd35438 & angle <= 16'd35455);
assign fi_addres[2055] = valid_point & (angle > 16'd35455 & angle <= 16'd35472);
assign fi_addres[2056] = valid_point & (angle > 16'd35472 & angle <= 16'd35489);
assign fi_addres[2057] = valid_point & (angle > 16'd35489 & angle <= 16'd35507);
assign fi_addres[2058] = valid_point & (angle > 16'd35507 & angle <= 16'd35525);
assign fi_addres[2059] = valid_point & (angle > 16'd35525 & angle <= 16'd35552);
assign fi_addres[2060] = valid_point & (angle > 16'd35552 & angle <= 16'd35570);
assign fi_addres[2061] = valid_point & (angle > 16'd35570 & angle <= 16'd35588);
assign fi_addres[2062] = valid_point & (angle > 16'd35588 & angle <= 16'd35606);
assign fi_addres[2063] = valid_point & (angle > 16'd35606 & angle <= 16'd35624);
assign fi_addres[2064] = valid_point & (angle > 16'd35624 & angle <= 16'd35642);
assign fi_addres[2065] = valid_point & (angle > 16'd35642 & angle <= 16'd35669);
assign fi_addres[2066] = valid_point & (angle > 16'd35669 & angle <= 16'd35687);
assign fi_addres[2067] = valid_point & (angle > 16'd35687 & angle <= 16'd35705);
assign fi_addres[2068] = valid_point & (angle > 16'd35705 & angle <= 16'd35723);
assign fi_addres[2069] = valid_point & (angle > 16'd35723 & angle <= 16'd35741);
assign fi_addres[2070] = valid_point & (angle > 16'd35741 & angle <= 16'd35771);
assign fi_addres[2071] = valid_point & (angle > 16'd35771 & angle <= 16'd35788);
assign fi_addres[2072] = valid_point & (angle > 16'd35788 & angle <= 16'd35804);
assign fi_addres[2073] = valid_point & (angle > 16'd35804 & angle <= 16'd35822);
assign fi_addres[2074] = valid_point & (angle > 16'd35822 & angle <= 16'd35840);
assign fi_addres[2075] = valid_point & (angle > 16'd35840 & angle <= 16'd35858);
assign fi_addres[2076] = valid_point & (angle > 16'd35858 & angle <= 16'd35876);
assign fi_addres[2077] = valid_point & (angle > 16'd35876 & angle <= 16'd35894);
assign fi_addres[2078] = valid_point & (angle > 16'd35894 & angle <= 16'd35924);
assign fi_addres[2079] = valid_point & (angle > 16'd35924 & angle <= 16'd35942);
assign fi_addres[2080] = valid_point & (angle > 16'd35942 & angle <= 16'd35975);
assign fi_addres[2081] = valid_point & (angle > 16'd35975 & angle <= 16'd36000);
        
endmodule
